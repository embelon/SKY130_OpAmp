magic
tech sky130A
magscale 1 2
timestamp 1695664993
<< error_p >>
rect -29 9233 29 9239
rect -29 9199 -17 9233
rect -29 9193 29 9199
rect -112 8052 112 8270
rect -29 7997 29 8003
rect -29 7963 -17 7997
rect -29 7957 29 7963
rect -112 6816 112 7034
rect -29 6761 29 6767
rect -29 6727 -17 6761
rect -29 6721 29 6727
rect -112 5580 112 5798
rect -29 5525 29 5531
rect -29 5491 -17 5525
rect -29 5485 29 5491
rect -112 4344 112 4562
rect -29 4289 29 4295
rect -29 4255 -17 4289
rect -29 4249 29 4255
rect -112 3108 112 3326
rect -29 3053 29 3059
rect -29 3019 -17 3053
rect -29 3013 29 3019
rect -112 1872 112 2090
rect -29 1817 29 1823
rect -29 1783 -17 1817
rect -29 1777 29 1783
rect -112 636 112 854
rect -29 581 29 587
rect -29 547 -17 581
rect -29 541 29 547
rect -112 -600 112 -382
rect -29 -655 29 -649
rect -29 -689 -17 -655
rect -29 -695 29 -689
rect -112 -1836 112 -1618
rect -29 -1891 29 -1885
rect -29 -1925 -17 -1891
rect -29 -1931 29 -1925
rect -112 -3072 112 -2854
rect -29 -3127 29 -3121
rect -29 -3161 -17 -3127
rect -29 -3167 29 -3161
rect -112 -4308 112 -4090
rect -29 -4363 29 -4357
rect -29 -4397 -17 -4363
rect -29 -4403 29 -4397
rect -112 -5544 112 -5326
rect -29 -5599 29 -5593
rect -29 -5633 -17 -5599
rect -29 -5639 29 -5633
rect -112 -6780 112 -6562
rect -29 -6835 29 -6829
rect -29 -6869 -17 -6835
rect -29 -6875 29 -6869
rect -112 -8016 112 -7798
rect -29 -8071 29 -8065
rect -29 -8105 -17 -8071
rect -29 -8111 29 -8105
rect -29 -9199 29 -9193
rect -29 -9233 -17 -9199
rect -29 -9239 29 -9233
<< nwell >>
rect -112 8052 112 9252
rect -112 6816 112 8016
rect -112 5580 112 6780
rect -112 4344 112 5544
rect -112 3108 112 4308
rect -112 1872 112 3072
rect -112 636 112 1836
rect -112 -600 112 600
rect -112 -1836 112 -636
rect -112 -3072 112 -1872
rect -112 -4308 112 -3108
rect -112 -5544 112 -4344
rect -112 -6780 112 -5580
rect -112 -8016 112 -6816
rect -112 -9252 112 -8052
<< pmos >>
rect -18 8152 18 9152
rect -18 6916 18 7916
rect -18 5680 18 6680
rect -18 4444 18 5444
rect -18 3208 18 4208
rect -18 1972 18 2972
rect -18 736 18 1736
rect -18 -500 18 500
rect -18 -1736 18 -736
rect -18 -2972 18 -1972
rect -18 -4208 18 -3208
rect -18 -5444 18 -4444
rect -18 -6680 18 -5680
rect -18 -7916 18 -6916
rect -18 -9152 18 -8152
<< pdiff >>
rect -76 9140 -18 9152
rect -76 8164 -64 9140
rect -30 8164 -18 9140
rect -76 8152 -18 8164
rect 18 9140 76 9152
rect 18 8164 30 9140
rect 64 8164 76 9140
rect 18 8152 76 8164
rect -76 7904 -18 7916
rect -76 6928 -64 7904
rect -30 6928 -18 7904
rect -76 6916 -18 6928
rect 18 7904 76 7916
rect 18 6928 30 7904
rect 64 6928 76 7904
rect 18 6916 76 6928
rect -76 6668 -18 6680
rect -76 5692 -64 6668
rect -30 5692 -18 6668
rect -76 5680 -18 5692
rect 18 6668 76 6680
rect 18 5692 30 6668
rect 64 5692 76 6668
rect 18 5680 76 5692
rect -76 5432 -18 5444
rect -76 4456 -64 5432
rect -30 4456 -18 5432
rect -76 4444 -18 4456
rect 18 5432 76 5444
rect 18 4456 30 5432
rect 64 4456 76 5432
rect 18 4444 76 4456
rect -76 4196 -18 4208
rect -76 3220 -64 4196
rect -30 3220 -18 4196
rect -76 3208 -18 3220
rect 18 4196 76 4208
rect 18 3220 30 4196
rect 64 3220 76 4196
rect 18 3208 76 3220
rect -76 2960 -18 2972
rect -76 1984 -64 2960
rect -30 1984 -18 2960
rect -76 1972 -18 1984
rect 18 2960 76 2972
rect 18 1984 30 2960
rect 64 1984 76 2960
rect 18 1972 76 1984
rect -76 1724 -18 1736
rect -76 748 -64 1724
rect -30 748 -18 1724
rect -76 736 -18 748
rect 18 1724 76 1736
rect 18 748 30 1724
rect 64 748 76 1724
rect 18 736 76 748
rect -76 488 -18 500
rect -76 -488 -64 488
rect -30 -488 -18 488
rect -76 -500 -18 -488
rect 18 488 76 500
rect 18 -488 30 488
rect 64 -488 76 488
rect 18 -500 76 -488
rect -76 -748 -18 -736
rect -76 -1724 -64 -748
rect -30 -1724 -18 -748
rect -76 -1736 -18 -1724
rect 18 -748 76 -736
rect 18 -1724 30 -748
rect 64 -1724 76 -748
rect 18 -1736 76 -1724
rect -76 -1984 -18 -1972
rect -76 -2960 -64 -1984
rect -30 -2960 -18 -1984
rect -76 -2972 -18 -2960
rect 18 -1984 76 -1972
rect 18 -2960 30 -1984
rect 64 -2960 76 -1984
rect 18 -2972 76 -2960
rect -76 -3220 -18 -3208
rect -76 -4196 -64 -3220
rect -30 -4196 -18 -3220
rect -76 -4208 -18 -4196
rect 18 -3220 76 -3208
rect 18 -4196 30 -3220
rect 64 -4196 76 -3220
rect 18 -4208 76 -4196
rect -76 -4456 -18 -4444
rect -76 -5432 -64 -4456
rect -30 -5432 -18 -4456
rect -76 -5444 -18 -5432
rect 18 -4456 76 -4444
rect 18 -5432 30 -4456
rect 64 -5432 76 -4456
rect 18 -5444 76 -5432
rect -76 -5692 -18 -5680
rect -76 -6668 -64 -5692
rect -30 -6668 -18 -5692
rect -76 -6680 -18 -6668
rect 18 -5692 76 -5680
rect 18 -6668 30 -5692
rect 64 -6668 76 -5692
rect 18 -6680 76 -6668
rect -76 -6928 -18 -6916
rect -76 -7904 -64 -6928
rect -30 -7904 -18 -6928
rect -76 -7916 -18 -7904
rect 18 -6928 76 -6916
rect 18 -7904 30 -6928
rect 64 -7904 76 -6928
rect 18 -7916 76 -7904
rect -76 -8164 -18 -8152
rect -76 -9140 -64 -8164
rect -30 -9140 -18 -8164
rect -76 -9152 -18 -9140
rect 18 -8164 76 -8152
rect 18 -9140 30 -8164
rect 64 -9140 76 -8164
rect 18 -9152 76 -9140
<< pdiffc >>
rect -64 8164 -30 9140
rect 30 8164 64 9140
rect -64 6928 -30 7904
rect 30 6928 64 7904
rect -64 5692 -30 6668
rect 30 5692 64 6668
rect -64 4456 -30 5432
rect 30 4456 64 5432
rect -64 3220 -30 4196
rect 30 3220 64 4196
rect -64 1984 -30 2960
rect 30 1984 64 2960
rect -64 748 -30 1724
rect 30 748 64 1724
rect -64 -488 -30 488
rect 30 -488 64 488
rect -64 -1724 -30 -748
rect 30 -1724 64 -748
rect -64 -2960 -30 -1984
rect 30 -2960 64 -1984
rect -64 -4196 -30 -3220
rect 30 -4196 64 -3220
rect -64 -5432 -30 -4456
rect 30 -5432 64 -4456
rect -64 -6668 -30 -5692
rect 30 -6668 64 -5692
rect -64 -7904 -30 -6928
rect 30 -7904 64 -6928
rect -64 -9140 -30 -8164
rect 30 -9140 64 -8164
<< poly >>
rect -33 9233 33 9249
rect -33 9199 -17 9233
rect 17 9199 33 9233
rect -33 9183 33 9199
rect -18 9152 18 9183
rect -18 8121 18 8152
rect -33 8105 33 8121
rect -33 8071 -17 8105
rect 17 8071 33 8105
rect -33 8055 33 8071
rect -33 7997 33 8013
rect -33 7963 -17 7997
rect 17 7963 33 7997
rect -33 7947 33 7963
rect -18 7916 18 7947
rect -18 6885 18 6916
rect -33 6869 33 6885
rect -33 6835 -17 6869
rect 17 6835 33 6869
rect -33 6819 33 6835
rect -33 6761 33 6777
rect -33 6727 -17 6761
rect 17 6727 33 6761
rect -33 6711 33 6727
rect -18 6680 18 6711
rect -18 5649 18 5680
rect -33 5633 33 5649
rect -33 5599 -17 5633
rect 17 5599 33 5633
rect -33 5583 33 5599
rect -33 5525 33 5541
rect -33 5491 -17 5525
rect 17 5491 33 5525
rect -33 5475 33 5491
rect -18 5444 18 5475
rect -18 4413 18 4444
rect -33 4397 33 4413
rect -33 4363 -17 4397
rect 17 4363 33 4397
rect -33 4347 33 4363
rect -33 4289 33 4305
rect -33 4255 -17 4289
rect 17 4255 33 4289
rect -33 4239 33 4255
rect -18 4208 18 4239
rect -18 3177 18 3208
rect -33 3161 33 3177
rect -33 3127 -17 3161
rect 17 3127 33 3161
rect -33 3111 33 3127
rect -33 3053 33 3069
rect -33 3019 -17 3053
rect 17 3019 33 3053
rect -33 3003 33 3019
rect -18 2972 18 3003
rect -18 1941 18 1972
rect -33 1925 33 1941
rect -33 1891 -17 1925
rect 17 1891 33 1925
rect -33 1875 33 1891
rect -33 1817 33 1833
rect -33 1783 -17 1817
rect 17 1783 33 1817
rect -33 1767 33 1783
rect -18 1736 18 1767
rect -18 705 18 736
rect -33 689 33 705
rect -33 655 -17 689
rect 17 655 33 689
rect -33 639 33 655
rect -33 581 33 597
rect -33 547 -17 581
rect 17 547 33 581
rect -33 531 33 547
rect -18 500 18 531
rect -18 -531 18 -500
rect -33 -547 33 -531
rect -33 -581 -17 -547
rect 17 -581 33 -547
rect -33 -597 33 -581
rect -33 -655 33 -639
rect -33 -689 -17 -655
rect 17 -689 33 -655
rect -33 -705 33 -689
rect -18 -736 18 -705
rect -18 -1767 18 -1736
rect -33 -1783 33 -1767
rect -33 -1817 -17 -1783
rect 17 -1817 33 -1783
rect -33 -1833 33 -1817
rect -33 -1891 33 -1875
rect -33 -1925 -17 -1891
rect 17 -1925 33 -1891
rect -33 -1941 33 -1925
rect -18 -1972 18 -1941
rect -18 -3003 18 -2972
rect -33 -3019 33 -3003
rect -33 -3053 -17 -3019
rect 17 -3053 33 -3019
rect -33 -3069 33 -3053
rect -33 -3127 33 -3111
rect -33 -3161 -17 -3127
rect 17 -3161 33 -3127
rect -33 -3177 33 -3161
rect -18 -3208 18 -3177
rect -18 -4239 18 -4208
rect -33 -4255 33 -4239
rect -33 -4289 -17 -4255
rect 17 -4289 33 -4255
rect -33 -4305 33 -4289
rect -33 -4363 33 -4347
rect -33 -4397 -17 -4363
rect 17 -4397 33 -4363
rect -33 -4413 33 -4397
rect -18 -4444 18 -4413
rect -18 -5475 18 -5444
rect -33 -5491 33 -5475
rect -33 -5525 -17 -5491
rect 17 -5525 33 -5491
rect -33 -5541 33 -5525
rect -33 -5599 33 -5583
rect -33 -5633 -17 -5599
rect 17 -5633 33 -5599
rect -33 -5649 33 -5633
rect -18 -5680 18 -5649
rect -18 -6711 18 -6680
rect -33 -6727 33 -6711
rect -33 -6761 -17 -6727
rect 17 -6761 33 -6727
rect -33 -6777 33 -6761
rect -33 -6835 33 -6819
rect -33 -6869 -17 -6835
rect 17 -6869 33 -6835
rect -33 -6885 33 -6869
rect -18 -6916 18 -6885
rect -18 -7947 18 -7916
rect -33 -7963 33 -7947
rect -33 -7997 -17 -7963
rect 17 -7997 33 -7963
rect -33 -8013 33 -7997
rect -33 -8071 33 -8055
rect -33 -8105 -17 -8071
rect 17 -8105 33 -8071
rect -33 -8121 33 -8105
rect -18 -8152 18 -8121
rect -18 -9183 18 -9152
rect -33 -9199 33 -9183
rect -33 -9233 -17 -9199
rect 17 -9233 33 -9199
rect -33 -9249 33 -9233
<< polycont >>
rect -17 9199 17 9233
rect -17 8071 17 8105
rect -17 7963 17 7997
rect -17 6835 17 6869
rect -17 6727 17 6761
rect -17 5599 17 5633
rect -17 5491 17 5525
rect -17 4363 17 4397
rect -17 4255 17 4289
rect -17 3127 17 3161
rect -17 3019 17 3053
rect -17 1891 17 1925
rect -17 1783 17 1817
rect -17 655 17 689
rect -17 547 17 581
rect -17 -581 17 -547
rect -17 -689 17 -655
rect -17 -1817 17 -1783
rect -17 -1925 17 -1891
rect -17 -3053 17 -3019
rect -17 -3161 17 -3127
rect -17 -4289 17 -4255
rect -17 -4397 17 -4363
rect -17 -5525 17 -5491
rect -17 -5633 17 -5599
rect -17 -6761 17 -6727
rect -17 -6869 17 -6835
rect -17 -7997 17 -7963
rect -17 -8105 17 -8071
rect -17 -9233 17 -9199
<< locali >>
rect -33 9199 -17 9233
rect 17 9199 33 9233
rect -64 9140 -30 9156
rect -64 8148 -30 8164
rect 30 9140 64 9156
rect 30 8148 64 8164
rect -33 8071 -17 8105
rect 17 8071 33 8105
rect -33 7963 -17 7997
rect 17 7963 33 7997
rect -64 7904 -30 7920
rect -64 6912 -30 6928
rect 30 7904 64 7920
rect 30 6912 64 6928
rect -33 6835 -17 6869
rect 17 6835 33 6869
rect -33 6727 -17 6761
rect 17 6727 33 6761
rect -64 6668 -30 6684
rect -64 5676 -30 5692
rect 30 6668 64 6684
rect 30 5676 64 5692
rect -33 5599 -17 5633
rect 17 5599 33 5633
rect -33 5491 -17 5525
rect 17 5491 33 5525
rect -64 5432 -30 5448
rect -64 4440 -30 4456
rect 30 5432 64 5448
rect 30 4440 64 4456
rect -33 4363 -17 4397
rect 17 4363 33 4397
rect -33 4255 -17 4289
rect 17 4255 33 4289
rect -64 4196 -30 4212
rect -64 3204 -30 3220
rect 30 4196 64 4212
rect 30 3204 64 3220
rect -33 3127 -17 3161
rect 17 3127 33 3161
rect -33 3019 -17 3053
rect 17 3019 33 3053
rect -64 2960 -30 2976
rect -64 1968 -30 1984
rect 30 2960 64 2976
rect 30 1968 64 1984
rect -33 1891 -17 1925
rect 17 1891 33 1925
rect -33 1783 -17 1817
rect 17 1783 33 1817
rect -64 1724 -30 1740
rect -64 732 -30 748
rect 30 1724 64 1740
rect 30 732 64 748
rect -33 655 -17 689
rect 17 655 33 689
rect -33 547 -17 581
rect 17 547 33 581
rect -64 488 -30 504
rect -64 -504 -30 -488
rect 30 488 64 504
rect 30 -504 64 -488
rect -33 -581 -17 -547
rect 17 -581 33 -547
rect -33 -689 -17 -655
rect 17 -689 33 -655
rect -64 -748 -30 -732
rect -64 -1740 -30 -1724
rect 30 -748 64 -732
rect 30 -1740 64 -1724
rect -33 -1817 -17 -1783
rect 17 -1817 33 -1783
rect -33 -1925 -17 -1891
rect 17 -1925 33 -1891
rect -64 -1984 -30 -1968
rect -64 -2976 -30 -2960
rect 30 -1984 64 -1968
rect 30 -2976 64 -2960
rect -33 -3053 -17 -3019
rect 17 -3053 33 -3019
rect -33 -3161 -17 -3127
rect 17 -3161 33 -3127
rect -64 -3220 -30 -3204
rect -64 -4212 -30 -4196
rect 30 -3220 64 -3204
rect 30 -4212 64 -4196
rect -33 -4289 -17 -4255
rect 17 -4289 33 -4255
rect -33 -4397 -17 -4363
rect 17 -4397 33 -4363
rect -64 -4456 -30 -4440
rect -64 -5448 -30 -5432
rect 30 -4456 64 -4440
rect 30 -5448 64 -5432
rect -33 -5525 -17 -5491
rect 17 -5525 33 -5491
rect -33 -5633 -17 -5599
rect 17 -5633 33 -5599
rect -64 -5692 -30 -5676
rect -64 -6684 -30 -6668
rect 30 -5692 64 -5676
rect 30 -6684 64 -6668
rect -33 -6761 -17 -6727
rect 17 -6761 33 -6727
rect -33 -6869 -17 -6835
rect 17 -6869 33 -6835
rect -64 -6928 -30 -6912
rect -64 -7920 -30 -7904
rect 30 -6928 64 -6912
rect 30 -7920 64 -7904
rect -33 -7997 -17 -7963
rect 17 -7997 33 -7963
rect -33 -8105 -17 -8071
rect 17 -8105 33 -8071
rect -64 -8164 -30 -8148
rect -64 -9156 -30 -9140
rect 30 -8164 64 -8148
rect 30 -9156 64 -9140
rect -33 -9233 -17 -9199
rect 17 -9233 33 -9199
<< viali >>
rect -17 9199 17 9233
rect -64 8164 -30 9140
rect 30 8164 64 9140
rect -17 8071 17 8105
rect -17 7963 17 7997
rect -64 6928 -30 7904
rect 30 6928 64 7904
rect -17 6835 17 6869
rect -17 6727 17 6761
rect -64 5692 -30 6668
rect 30 5692 64 6668
rect -17 5599 17 5633
rect -17 5491 17 5525
rect -64 4456 -30 5432
rect 30 4456 64 5432
rect -17 4363 17 4397
rect -17 4255 17 4289
rect -64 3220 -30 4196
rect 30 3220 64 4196
rect -17 3127 17 3161
rect -17 3019 17 3053
rect -64 1984 -30 2960
rect 30 1984 64 2960
rect -17 1891 17 1925
rect -17 1783 17 1817
rect -64 748 -30 1724
rect 30 748 64 1724
rect -17 655 17 689
rect -17 547 17 581
rect -64 -488 -30 488
rect 30 -488 64 488
rect -17 -581 17 -547
rect -17 -689 17 -655
rect -64 -1724 -30 -748
rect 30 -1724 64 -748
rect -17 -1817 17 -1783
rect -17 -1925 17 -1891
rect -64 -2960 -30 -1984
rect 30 -2960 64 -1984
rect -17 -3053 17 -3019
rect -17 -3161 17 -3127
rect -64 -4196 -30 -3220
rect 30 -4196 64 -3220
rect -17 -4289 17 -4255
rect -17 -4397 17 -4363
rect -64 -5432 -30 -4456
rect 30 -5432 64 -4456
rect -17 -5525 17 -5491
rect -17 -5633 17 -5599
rect -64 -6668 -30 -5692
rect 30 -6668 64 -5692
rect -17 -6761 17 -6727
rect -17 -6869 17 -6835
rect -64 -7904 -30 -6928
rect 30 -7904 64 -6928
rect -17 -7997 17 -7963
rect -17 -8105 17 -8071
rect -64 -9140 -30 -8164
rect 30 -9140 64 -8164
rect -17 -9233 17 -9199
<< metal1 >>
rect -29 9233 29 9239
rect -29 9199 -17 9233
rect 17 9199 29 9233
rect -29 9193 29 9199
rect -70 9140 -24 9152
rect -70 8164 -64 9140
rect -30 8164 -24 9140
rect -70 8152 -24 8164
rect 24 9140 70 9152
rect 24 8164 30 9140
rect 64 8164 70 9140
rect 24 8152 70 8164
rect -29 8105 29 8111
rect -29 8071 -17 8105
rect 17 8071 29 8105
rect -29 8065 29 8071
rect -29 7997 29 8003
rect -29 7963 -17 7997
rect 17 7963 29 7997
rect -29 7957 29 7963
rect -70 7904 -24 7916
rect -70 6928 -64 7904
rect -30 6928 -24 7904
rect -70 6916 -24 6928
rect 24 7904 70 7916
rect 24 6928 30 7904
rect 64 6928 70 7904
rect 24 6916 70 6928
rect -29 6869 29 6875
rect -29 6835 -17 6869
rect 17 6835 29 6869
rect -29 6829 29 6835
rect -29 6761 29 6767
rect -29 6727 -17 6761
rect 17 6727 29 6761
rect -29 6721 29 6727
rect -70 6668 -24 6680
rect -70 5692 -64 6668
rect -30 5692 -24 6668
rect -70 5680 -24 5692
rect 24 6668 70 6680
rect 24 5692 30 6668
rect 64 5692 70 6668
rect 24 5680 70 5692
rect -29 5633 29 5639
rect -29 5599 -17 5633
rect 17 5599 29 5633
rect -29 5593 29 5599
rect -29 5525 29 5531
rect -29 5491 -17 5525
rect 17 5491 29 5525
rect -29 5485 29 5491
rect -70 5432 -24 5444
rect -70 4456 -64 5432
rect -30 4456 -24 5432
rect -70 4444 -24 4456
rect 24 5432 70 5444
rect 24 4456 30 5432
rect 64 4456 70 5432
rect 24 4444 70 4456
rect -29 4397 29 4403
rect -29 4363 -17 4397
rect 17 4363 29 4397
rect -29 4357 29 4363
rect -29 4289 29 4295
rect -29 4255 -17 4289
rect 17 4255 29 4289
rect -29 4249 29 4255
rect -70 4196 -24 4208
rect -70 3220 -64 4196
rect -30 3220 -24 4196
rect -70 3208 -24 3220
rect 24 4196 70 4208
rect 24 3220 30 4196
rect 64 3220 70 4196
rect 24 3208 70 3220
rect -29 3161 29 3167
rect -29 3127 -17 3161
rect 17 3127 29 3161
rect -29 3121 29 3127
rect -29 3053 29 3059
rect -29 3019 -17 3053
rect 17 3019 29 3053
rect -29 3013 29 3019
rect -70 2960 -24 2972
rect -70 1984 -64 2960
rect -30 1984 -24 2960
rect -70 1972 -24 1984
rect 24 2960 70 2972
rect 24 1984 30 2960
rect 64 1984 70 2960
rect 24 1972 70 1984
rect -29 1925 29 1931
rect -29 1891 -17 1925
rect 17 1891 29 1925
rect -29 1885 29 1891
rect -29 1817 29 1823
rect -29 1783 -17 1817
rect 17 1783 29 1817
rect -29 1777 29 1783
rect -70 1724 -24 1736
rect -70 748 -64 1724
rect -30 748 -24 1724
rect -70 736 -24 748
rect 24 1724 70 1736
rect 24 748 30 1724
rect 64 748 70 1724
rect 24 736 70 748
rect -29 689 29 695
rect -29 655 -17 689
rect 17 655 29 689
rect -29 649 29 655
rect -29 581 29 587
rect -29 547 -17 581
rect 17 547 29 581
rect -29 541 29 547
rect -70 488 -24 500
rect -70 -488 -64 488
rect -30 -488 -24 488
rect -70 -500 -24 -488
rect 24 488 70 500
rect 24 -488 30 488
rect 64 -488 70 488
rect 24 -500 70 -488
rect -29 -547 29 -541
rect -29 -581 -17 -547
rect 17 -581 29 -547
rect -29 -587 29 -581
rect -29 -655 29 -649
rect -29 -689 -17 -655
rect 17 -689 29 -655
rect -29 -695 29 -689
rect -70 -748 -24 -736
rect -70 -1724 -64 -748
rect -30 -1724 -24 -748
rect -70 -1736 -24 -1724
rect 24 -748 70 -736
rect 24 -1724 30 -748
rect 64 -1724 70 -748
rect 24 -1736 70 -1724
rect -29 -1783 29 -1777
rect -29 -1817 -17 -1783
rect 17 -1817 29 -1783
rect -29 -1823 29 -1817
rect -29 -1891 29 -1885
rect -29 -1925 -17 -1891
rect 17 -1925 29 -1891
rect -29 -1931 29 -1925
rect -70 -1984 -24 -1972
rect -70 -2960 -64 -1984
rect -30 -2960 -24 -1984
rect -70 -2972 -24 -2960
rect 24 -1984 70 -1972
rect 24 -2960 30 -1984
rect 64 -2960 70 -1984
rect 24 -2972 70 -2960
rect -29 -3019 29 -3013
rect -29 -3053 -17 -3019
rect 17 -3053 29 -3019
rect -29 -3059 29 -3053
rect -29 -3127 29 -3121
rect -29 -3161 -17 -3127
rect 17 -3161 29 -3127
rect -29 -3167 29 -3161
rect -70 -3220 -24 -3208
rect -70 -4196 -64 -3220
rect -30 -4196 -24 -3220
rect -70 -4208 -24 -4196
rect 24 -3220 70 -3208
rect 24 -4196 30 -3220
rect 64 -4196 70 -3220
rect 24 -4208 70 -4196
rect -29 -4255 29 -4249
rect -29 -4289 -17 -4255
rect 17 -4289 29 -4255
rect -29 -4295 29 -4289
rect -29 -4363 29 -4357
rect -29 -4397 -17 -4363
rect 17 -4397 29 -4363
rect -29 -4403 29 -4397
rect -70 -4456 -24 -4444
rect -70 -5432 -64 -4456
rect -30 -5432 -24 -4456
rect -70 -5444 -24 -5432
rect 24 -4456 70 -4444
rect 24 -5432 30 -4456
rect 64 -5432 70 -4456
rect 24 -5444 70 -5432
rect -29 -5491 29 -5485
rect -29 -5525 -17 -5491
rect 17 -5525 29 -5491
rect -29 -5531 29 -5525
rect -29 -5599 29 -5593
rect -29 -5633 -17 -5599
rect 17 -5633 29 -5599
rect -29 -5639 29 -5633
rect -70 -5692 -24 -5680
rect -70 -6668 -64 -5692
rect -30 -6668 -24 -5692
rect -70 -6680 -24 -6668
rect 24 -5692 70 -5680
rect 24 -6668 30 -5692
rect 64 -6668 70 -5692
rect 24 -6680 70 -6668
rect -29 -6727 29 -6721
rect -29 -6761 -17 -6727
rect 17 -6761 29 -6727
rect -29 -6767 29 -6761
rect -29 -6835 29 -6829
rect -29 -6869 -17 -6835
rect 17 -6869 29 -6835
rect -29 -6875 29 -6869
rect -70 -6928 -24 -6916
rect -70 -7904 -64 -6928
rect -30 -7904 -24 -6928
rect -70 -7916 -24 -7904
rect 24 -6928 70 -6916
rect 24 -7904 30 -6928
rect 64 -7904 70 -6928
rect 24 -7916 70 -7904
rect -29 -7963 29 -7957
rect -29 -7997 -17 -7963
rect 17 -7997 29 -7963
rect -29 -8003 29 -7997
rect -29 -8071 29 -8065
rect -29 -8105 -17 -8071
rect 17 -8105 29 -8071
rect -29 -8111 29 -8105
rect -70 -8164 -24 -8152
rect -70 -9140 -64 -8164
rect -30 -9140 -24 -8164
rect -70 -9152 -24 -9140
rect 24 -8164 70 -8152
rect 24 -9140 30 -8164
rect 64 -9140 70 -8164
rect 24 -9152 70 -9140
rect -29 -9199 29 -9193
rect -29 -9233 -17 -9199
rect 17 -9233 29 -9199
rect -29 -9239 29 -9233
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 5.0 l 0.18 m 15 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
