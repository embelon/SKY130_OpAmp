VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO opamp_cascode
  CLASS BLOCK ;
  FOREIGN opamp_cascode ;
  ORIGIN -164.000 -70.000 ;
  SIZE 366.000 BY 655.000 ;
  PIN IN_P
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 64.799995 ;
    PORT
      LAYER met3 ;
        RECT 164.000 70.000 174.000 80.000 ;
    END
  END IN_P
  PIN IN_M
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 27.000000 ;
    PORT
      LAYER met3 ;
        RECT 164.000 90.000 174.000 100.000 ;
    END
  END IN_M
  PIN VCC
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 164.000 695.000 191.000 705.000 ;
    END
  END VCC
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 164.000 715.000 273.000 725.000 ;
    END
  END VSS
  PIN OUT
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 87.000000 ;
    PORT
      LAYER met3 ;
        RECT 164.000 450.000 174.000 460.000 ;
    END
  END OUT
  PIN VB_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2550.000000 ;
    PORT
      LAYER met3 ;
        RECT 164.000 430.000 174.000 440.000 ;
    END
  END VB_A
  PIN VB_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2550.000000 ;
    PORT
      LAYER met3 ;
        RECT 164.000 560.000 174.000 570.000 ;
    END
  END VB_B
  PIN IB
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 450.000000 ;
    ANTENNADIFFAREA 5.800000 ;
    PORT
      LAYER met3 ;
        RECT 164.000 270.000 174.000 280.000 ;
    END
  END IB
  OBS
      LAYER li1 ;
        RECT 201.500 79.095 523.700 719.400 ;
      LAYER met1 ;
        RECT 201.950 74.500 524.500 722.000 ;
      LAYER met2 ;
        RECT 180.000 71.950 524.000 725.000 ;
      LAYER met3 ;
        RECT 174.000 705.400 273.050 714.600 ;
        RECT 191.400 694.600 273.050 705.400 ;
        RECT 174.000 570.400 273.050 694.600 ;
        RECT 174.400 559.600 273.050 570.400 ;
        RECT 174.000 460.400 273.050 559.600 ;
        RECT 174.400 449.600 273.050 460.400 ;
        RECT 174.000 440.400 273.050 449.600 ;
        RECT 174.400 429.600 273.050 440.400 ;
        RECT 174.000 280.400 273.050 429.600 ;
        RECT 174.400 269.600 273.050 280.400 ;
        RECT 174.000 100.400 273.050 269.600 ;
        RECT 174.400 89.600 273.050 100.400 ;
        RECT 174.000 80.400 273.050 89.600 ;
        RECT 174.400 70.000 273.050 80.400 ;
  END
END opamp_cascode
END LIBRARY

