** sch_path: ../opamp_cascode_ac_openloop.sch
**.subckt opamp_cascode_ac_openloop
C1 Vout GND 1p m=1
V1 Vfb Vm 0 AC 1
.save i(v1)
R1 Vfb Vout 100k m=1
R2 Vp Vfb 100k m=1
I0 IBIAS GND 45u
x1 Vp Vm VCC GND Vout VB_A VB_B IBIAS opamp_cascode
**** begin user architecture code


Vsupply VCC GND 1.8
VbiasA VB_A GND 0.2
VbiasB VB_B GND 1.1
Vin Vp GND 0.9
.include ../opamp_cascode.spice
.control
  save all
  ac dec 10 1 1G
  let T = v(Vfb) / v(Vm)
  let mag = db(T)
  let phase = 180*cph(T)/pi
  plot mag phase xlog
  meas ac margin find phase when mag=0
  meas ac GBW when mag=0
.endc



.param mc_mm_switch=1
.param mc_pr_switch=0
.include ~/.volare/sky130A/libs.tech/ngspice/corners/tt.spice
.include ~/.volare/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include ~/.volare/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include ~/.volare/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice

**** end user architecture code
**.ends
.GLOBAL GND
.end
