magic
tech sky130A
magscale 1 2
timestamp 1695661682
<< nwell >>
rect -696 -9371 696 9371
<< pmos >>
rect -500 8152 500 9152
rect -500 6916 500 7916
rect -500 5680 500 6680
rect -500 4444 500 5444
rect -500 3208 500 4208
rect -500 1972 500 2972
rect -500 736 500 1736
rect -500 -500 500 500
rect -500 -1736 500 -736
rect -500 -2972 500 -1972
rect -500 -4208 500 -3208
rect -500 -5444 500 -4444
rect -500 -6680 500 -5680
rect -500 -7916 500 -6916
rect -500 -9152 500 -8152
<< pdiff >>
rect -558 9140 -500 9152
rect -558 8164 -546 9140
rect -512 8164 -500 9140
rect -558 8152 -500 8164
rect 500 9140 558 9152
rect 500 8164 512 9140
rect 546 8164 558 9140
rect 500 8152 558 8164
rect -558 7904 -500 7916
rect -558 6928 -546 7904
rect -512 6928 -500 7904
rect -558 6916 -500 6928
rect 500 7904 558 7916
rect 500 6928 512 7904
rect 546 6928 558 7904
rect 500 6916 558 6928
rect -558 6668 -500 6680
rect -558 5692 -546 6668
rect -512 5692 -500 6668
rect -558 5680 -500 5692
rect 500 6668 558 6680
rect 500 5692 512 6668
rect 546 5692 558 6668
rect 500 5680 558 5692
rect -558 5432 -500 5444
rect -558 4456 -546 5432
rect -512 4456 -500 5432
rect -558 4444 -500 4456
rect 500 5432 558 5444
rect 500 4456 512 5432
rect 546 4456 558 5432
rect 500 4444 558 4456
rect -558 4196 -500 4208
rect -558 3220 -546 4196
rect -512 3220 -500 4196
rect -558 3208 -500 3220
rect 500 4196 558 4208
rect 500 3220 512 4196
rect 546 3220 558 4196
rect 500 3208 558 3220
rect -558 2960 -500 2972
rect -558 1984 -546 2960
rect -512 1984 -500 2960
rect -558 1972 -500 1984
rect 500 2960 558 2972
rect 500 1984 512 2960
rect 546 1984 558 2960
rect 500 1972 558 1984
rect -558 1724 -500 1736
rect -558 748 -546 1724
rect -512 748 -500 1724
rect -558 736 -500 748
rect 500 1724 558 1736
rect 500 748 512 1724
rect 546 748 558 1724
rect 500 736 558 748
rect -558 488 -500 500
rect -558 -488 -546 488
rect -512 -488 -500 488
rect -558 -500 -500 -488
rect 500 488 558 500
rect 500 -488 512 488
rect 546 -488 558 488
rect 500 -500 558 -488
rect -558 -748 -500 -736
rect -558 -1724 -546 -748
rect -512 -1724 -500 -748
rect -558 -1736 -500 -1724
rect 500 -748 558 -736
rect 500 -1724 512 -748
rect 546 -1724 558 -748
rect 500 -1736 558 -1724
rect -558 -1984 -500 -1972
rect -558 -2960 -546 -1984
rect -512 -2960 -500 -1984
rect -558 -2972 -500 -2960
rect 500 -1984 558 -1972
rect 500 -2960 512 -1984
rect 546 -2960 558 -1984
rect 500 -2972 558 -2960
rect -558 -3220 -500 -3208
rect -558 -4196 -546 -3220
rect -512 -4196 -500 -3220
rect -558 -4208 -500 -4196
rect 500 -3220 558 -3208
rect 500 -4196 512 -3220
rect 546 -4196 558 -3220
rect 500 -4208 558 -4196
rect -558 -4456 -500 -4444
rect -558 -5432 -546 -4456
rect -512 -5432 -500 -4456
rect -558 -5444 -500 -5432
rect 500 -4456 558 -4444
rect 500 -5432 512 -4456
rect 546 -5432 558 -4456
rect 500 -5444 558 -5432
rect -558 -5692 -500 -5680
rect -558 -6668 -546 -5692
rect -512 -6668 -500 -5692
rect -558 -6680 -500 -6668
rect 500 -5692 558 -5680
rect 500 -6668 512 -5692
rect 546 -6668 558 -5692
rect 500 -6680 558 -6668
rect -558 -6928 -500 -6916
rect -558 -7904 -546 -6928
rect -512 -7904 -500 -6928
rect -558 -7916 -500 -7904
rect 500 -6928 558 -6916
rect 500 -7904 512 -6928
rect 546 -7904 558 -6928
rect 500 -7916 558 -7904
rect -558 -8164 -500 -8152
rect -558 -9140 -546 -8164
rect -512 -9140 -500 -8164
rect -558 -9152 -500 -9140
rect 500 -8164 558 -8152
rect 500 -9140 512 -8164
rect 546 -9140 558 -8164
rect 500 -9152 558 -9140
<< pdiffc >>
rect -546 8164 -512 9140
rect 512 8164 546 9140
rect -546 6928 -512 7904
rect 512 6928 546 7904
rect -546 5692 -512 6668
rect 512 5692 546 6668
rect -546 4456 -512 5432
rect 512 4456 546 5432
rect -546 3220 -512 4196
rect 512 3220 546 4196
rect -546 1984 -512 2960
rect 512 1984 546 2960
rect -546 748 -512 1724
rect 512 748 546 1724
rect -546 -488 -512 488
rect 512 -488 546 488
rect -546 -1724 -512 -748
rect 512 -1724 546 -748
rect -546 -2960 -512 -1984
rect 512 -2960 546 -1984
rect -546 -4196 -512 -3220
rect 512 -4196 546 -3220
rect -546 -5432 -512 -4456
rect 512 -5432 546 -4456
rect -546 -6668 -512 -5692
rect 512 -6668 546 -5692
rect -546 -7904 -512 -6928
rect 512 -7904 546 -6928
rect -546 -9140 -512 -8164
rect 512 -9140 546 -8164
<< nsubdiff >>
rect -660 9301 -564 9335
rect 564 9301 660 9335
rect -660 9239 -626 9301
rect 626 9239 660 9301
rect -660 -9301 -626 -9239
rect 626 -9301 660 -9239
rect -660 -9335 -564 -9301
rect 564 -9335 660 -9301
<< nsubdiffcont >>
rect -564 9301 564 9335
rect -660 -9239 -626 9239
rect 626 -9239 660 9239
rect -564 -9335 564 -9301
<< poly >>
rect -500 9233 500 9249
rect -500 9199 -484 9233
rect 484 9199 500 9233
rect -500 9152 500 9199
rect -500 8105 500 8152
rect -500 8071 -484 8105
rect 484 8071 500 8105
rect -500 8055 500 8071
rect -500 7997 500 8013
rect -500 7963 -484 7997
rect 484 7963 500 7997
rect -500 7916 500 7963
rect -500 6869 500 6916
rect -500 6835 -484 6869
rect 484 6835 500 6869
rect -500 6819 500 6835
rect -500 6761 500 6777
rect -500 6727 -484 6761
rect 484 6727 500 6761
rect -500 6680 500 6727
rect -500 5633 500 5680
rect -500 5599 -484 5633
rect 484 5599 500 5633
rect -500 5583 500 5599
rect -500 5525 500 5541
rect -500 5491 -484 5525
rect 484 5491 500 5525
rect -500 5444 500 5491
rect -500 4397 500 4444
rect -500 4363 -484 4397
rect 484 4363 500 4397
rect -500 4347 500 4363
rect -500 4289 500 4305
rect -500 4255 -484 4289
rect 484 4255 500 4289
rect -500 4208 500 4255
rect -500 3161 500 3208
rect -500 3127 -484 3161
rect 484 3127 500 3161
rect -500 3111 500 3127
rect -500 3053 500 3069
rect -500 3019 -484 3053
rect 484 3019 500 3053
rect -500 2972 500 3019
rect -500 1925 500 1972
rect -500 1891 -484 1925
rect 484 1891 500 1925
rect -500 1875 500 1891
rect -500 1817 500 1833
rect -500 1783 -484 1817
rect 484 1783 500 1817
rect -500 1736 500 1783
rect -500 689 500 736
rect -500 655 -484 689
rect 484 655 500 689
rect -500 639 500 655
rect -500 581 500 597
rect -500 547 -484 581
rect 484 547 500 581
rect -500 500 500 547
rect -500 -547 500 -500
rect -500 -581 -484 -547
rect 484 -581 500 -547
rect -500 -597 500 -581
rect -500 -655 500 -639
rect -500 -689 -484 -655
rect 484 -689 500 -655
rect -500 -736 500 -689
rect -500 -1783 500 -1736
rect -500 -1817 -484 -1783
rect 484 -1817 500 -1783
rect -500 -1833 500 -1817
rect -500 -1891 500 -1875
rect -500 -1925 -484 -1891
rect 484 -1925 500 -1891
rect -500 -1972 500 -1925
rect -500 -3019 500 -2972
rect -500 -3053 -484 -3019
rect 484 -3053 500 -3019
rect -500 -3069 500 -3053
rect -500 -3127 500 -3111
rect -500 -3161 -484 -3127
rect 484 -3161 500 -3127
rect -500 -3208 500 -3161
rect -500 -4255 500 -4208
rect -500 -4289 -484 -4255
rect 484 -4289 500 -4255
rect -500 -4305 500 -4289
rect -500 -4363 500 -4347
rect -500 -4397 -484 -4363
rect 484 -4397 500 -4363
rect -500 -4444 500 -4397
rect -500 -5491 500 -5444
rect -500 -5525 -484 -5491
rect 484 -5525 500 -5491
rect -500 -5541 500 -5525
rect -500 -5599 500 -5583
rect -500 -5633 -484 -5599
rect 484 -5633 500 -5599
rect -500 -5680 500 -5633
rect -500 -6727 500 -6680
rect -500 -6761 -484 -6727
rect 484 -6761 500 -6727
rect -500 -6777 500 -6761
rect -500 -6835 500 -6819
rect -500 -6869 -484 -6835
rect 484 -6869 500 -6835
rect -500 -6916 500 -6869
rect -500 -7963 500 -7916
rect -500 -7997 -484 -7963
rect 484 -7997 500 -7963
rect -500 -8013 500 -7997
rect -500 -8071 500 -8055
rect -500 -8105 -484 -8071
rect 484 -8105 500 -8071
rect -500 -8152 500 -8105
rect -500 -9199 500 -9152
rect -500 -9233 -484 -9199
rect 484 -9233 500 -9199
rect -500 -9249 500 -9233
<< polycont >>
rect -484 9199 484 9233
rect -484 8071 484 8105
rect -484 7963 484 7997
rect -484 6835 484 6869
rect -484 6727 484 6761
rect -484 5599 484 5633
rect -484 5491 484 5525
rect -484 4363 484 4397
rect -484 4255 484 4289
rect -484 3127 484 3161
rect -484 3019 484 3053
rect -484 1891 484 1925
rect -484 1783 484 1817
rect -484 655 484 689
rect -484 547 484 581
rect -484 -581 484 -547
rect -484 -689 484 -655
rect -484 -1817 484 -1783
rect -484 -1925 484 -1891
rect -484 -3053 484 -3019
rect -484 -3161 484 -3127
rect -484 -4289 484 -4255
rect -484 -4397 484 -4363
rect -484 -5525 484 -5491
rect -484 -5633 484 -5599
rect -484 -6761 484 -6727
rect -484 -6869 484 -6835
rect -484 -7997 484 -7963
rect -484 -8105 484 -8071
rect -484 -9233 484 -9199
<< locali >>
rect -660 9301 -564 9335
rect 564 9301 660 9335
rect -660 9239 -626 9301
rect 626 9239 660 9301
rect -500 9199 -484 9233
rect 484 9199 500 9233
rect -546 9140 -512 9156
rect -546 8148 -512 8164
rect 512 9140 546 9156
rect 512 8148 546 8164
rect -500 8071 -484 8105
rect 484 8071 500 8105
rect -500 7963 -484 7997
rect 484 7963 500 7997
rect -546 7904 -512 7920
rect -546 6912 -512 6928
rect 512 7904 546 7920
rect 512 6912 546 6928
rect -500 6835 -484 6869
rect 484 6835 500 6869
rect -500 6727 -484 6761
rect 484 6727 500 6761
rect -546 6668 -512 6684
rect -546 5676 -512 5692
rect 512 6668 546 6684
rect 512 5676 546 5692
rect -500 5599 -484 5633
rect 484 5599 500 5633
rect -500 5491 -484 5525
rect 484 5491 500 5525
rect -546 5432 -512 5448
rect -546 4440 -512 4456
rect 512 5432 546 5448
rect 512 4440 546 4456
rect -500 4363 -484 4397
rect 484 4363 500 4397
rect -500 4255 -484 4289
rect 484 4255 500 4289
rect -546 4196 -512 4212
rect -546 3204 -512 3220
rect 512 4196 546 4212
rect 512 3204 546 3220
rect -500 3127 -484 3161
rect 484 3127 500 3161
rect -500 3019 -484 3053
rect 484 3019 500 3053
rect -546 2960 -512 2976
rect -546 1968 -512 1984
rect 512 2960 546 2976
rect 512 1968 546 1984
rect -500 1891 -484 1925
rect 484 1891 500 1925
rect -500 1783 -484 1817
rect 484 1783 500 1817
rect -546 1724 -512 1740
rect -546 732 -512 748
rect 512 1724 546 1740
rect 512 732 546 748
rect -500 655 -484 689
rect 484 655 500 689
rect -500 547 -484 581
rect 484 547 500 581
rect -546 488 -512 504
rect -546 -504 -512 -488
rect 512 488 546 504
rect 512 -504 546 -488
rect -500 -581 -484 -547
rect 484 -581 500 -547
rect -500 -689 -484 -655
rect 484 -689 500 -655
rect -546 -748 -512 -732
rect -546 -1740 -512 -1724
rect 512 -748 546 -732
rect 512 -1740 546 -1724
rect -500 -1817 -484 -1783
rect 484 -1817 500 -1783
rect -500 -1925 -484 -1891
rect 484 -1925 500 -1891
rect -546 -1984 -512 -1968
rect -546 -2976 -512 -2960
rect 512 -1984 546 -1968
rect 512 -2976 546 -2960
rect -500 -3053 -484 -3019
rect 484 -3053 500 -3019
rect -500 -3161 -484 -3127
rect 484 -3161 500 -3127
rect -546 -3220 -512 -3204
rect -546 -4212 -512 -4196
rect 512 -3220 546 -3204
rect 512 -4212 546 -4196
rect -500 -4289 -484 -4255
rect 484 -4289 500 -4255
rect -500 -4397 -484 -4363
rect 484 -4397 500 -4363
rect -546 -4456 -512 -4440
rect -546 -5448 -512 -5432
rect 512 -4456 546 -4440
rect 512 -5448 546 -5432
rect -500 -5525 -484 -5491
rect 484 -5525 500 -5491
rect -500 -5633 -484 -5599
rect 484 -5633 500 -5599
rect -546 -5692 -512 -5676
rect -546 -6684 -512 -6668
rect 512 -5692 546 -5676
rect 512 -6684 546 -6668
rect -500 -6761 -484 -6727
rect 484 -6761 500 -6727
rect -500 -6869 -484 -6835
rect 484 -6869 500 -6835
rect -546 -6928 -512 -6912
rect -546 -7920 -512 -7904
rect 512 -6928 546 -6912
rect 512 -7920 546 -7904
rect -500 -7997 -484 -7963
rect 484 -7997 500 -7963
rect -500 -8105 -484 -8071
rect 484 -8105 500 -8071
rect -546 -8164 -512 -8148
rect -546 -9156 -512 -9140
rect 512 -8164 546 -8148
rect 512 -9156 546 -9140
rect -500 -9233 -484 -9199
rect 484 -9233 500 -9199
rect -660 -9301 -626 -9239
rect 626 -9301 660 -9239
rect -660 -9335 -564 -9301
rect 564 -9335 660 -9301
<< viali >>
rect -484 9199 484 9233
rect -546 8164 -512 9140
rect 512 8164 546 9140
rect -484 8071 484 8105
rect -484 7963 484 7997
rect -546 6928 -512 7904
rect 512 6928 546 7904
rect -484 6835 484 6869
rect -484 6727 484 6761
rect -546 5692 -512 6668
rect 512 5692 546 6668
rect -484 5599 484 5633
rect -484 5491 484 5525
rect -546 4456 -512 5432
rect 512 4456 546 5432
rect -484 4363 484 4397
rect -484 4255 484 4289
rect -546 3220 -512 4196
rect 512 3220 546 4196
rect -484 3127 484 3161
rect -484 3019 484 3053
rect -546 1984 -512 2960
rect 512 1984 546 2960
rect -484 1891 484 1925
rect -484 1783 484 1817
rect -546 748 -512 1724
rect 512 748 546 1724
rect -484 655 484 689
rect -484 547 484 581
rect -546 -488 -512 488
rect 512 -488 546 488
rect -484 -581 484 -547
rect -484 -689 484 -655
rect -546 -1724 -512 -748
rect 512 -1724 546 -748
rect -484 -1817 484 -1783
rect -484 -1925 484 -1891
rect -546 -2960 -512 -1984
rect 512 -2960 546 -1984
rect -484 -3053 484 -3019
rect -484 -3161 484 -3127
rect -546 -4196 -512 -3220
rect 512 -4196 546 -3220
rect -484 -4289 484 -4255
rect -484 -4397 484 -4363
rect -546 -5432 -512 -4456
rect 512 -5432 546 -4456
rect -484 -5525 484 -5491
rect -484 -5633 484 -5599
rect -546 -6668 -512 -5692
rect 512 -6668 546 -5692
rect -484 -6761 484 -6727
rect -484 -6869 484 -6835
rect -546 -7904 -512 -6928
rect 512 -7904 546 -6928
rect -484 -7997 484 -7963
rect -484 -8105 484 -8071
rect -546 -9140 -512 -8164
rect 512 -9140 546 -8164
rect -484 -9233 484 -9199
<< metal1 >>
rect -496 9233 496 9239
rect -496 9199 -484 9233
rect 484 9199 496 9233
rect -496 9193 496 9199
rect -552 9140 -506 9152
rect -552 8164 -546 9140
rect -512 8164 -506 9140
rect -552 8152 -506 8164
rect 506 9140 552 9152
rect 506 8164 512 9140
rect 546 8164 552 9140
rect 506 8152 552 8164
rect -496 8105 496 8111
rect -496 8071 -484 8105
rect 484 8071 496 8105
rect -496 8065 496 8071
rect -496 7997 496 8003
rect -496 7963 -484 7997
rect 484 7963 496 7997
rect -496 7957 496 7963
rect -552 7904 -506 7916
rect -552 6928 -546 7904
rect -512 6928 -506 7904
rect -552 6916 -506 6928
rect 506 7904 552 7916
rect 506 6928 512 7904
rect 546 6928 552 7904
rect 506 6916 552 6928
rect -496 6869 496 6875
rect -496 6835 -484 6869
rect 484 6835 496 6869
rect -496 6829 496 6835
rect -496 6761 496 6767
rect -496 6727 -484 6761
rect 484 6727 496 6761
rect -496 6721 496 6727
rect -552 6668 -506 6680
rect -552 5692 -546 6668
rect -512 5692 -506 6668
rect -552 5680 -506 5692
rect 506 6668 552 6680
rect 506 5692 512 6668
rect 546 5692 552 6668
rect 506 5680 552 5692
rect -496 5633 496 5639
rect -496 5599 -484 5633
rect 484 5599 496 5633
rect -496 5593 496 5599
rect -496 5525 496 5531
rect -496 5491 -484 5525
rect 484 5491 496 5525
rect -496 5485 496 5491
rect -552 5432 -506 5444
rect -552 4456 -546 5432
rect -512 4456 -506 5432
rect -552 4444 -506 4456
rect 506 5432 552 5444
rect 506 4456 512 5432
rect 546 4456 552 5432
rect 506 4444 552 4456
rect -496 4397 496 4403
rect -496 4363 -484 4397
rect 484 4363 496 4397
rect -496 4357 496 4363
rect -496 4289 496 4295
rect -496 4255 -484 4289
rect 484 4255 496 4289
rect -496 4249 496 4255
rect -552 4196 -506 4208
rect -552 3220 -546 4196
rect -512 3220 -506 4196
rect -552 3208 -506 3220
rect 506 4196 552 4208
rect 506 3220 512 4196
rect 546 3220 552 4196
rect 506 3208 552 3220
rect -496 3161 496 3167
rect -496 3127 -484 3161
rect 484 3127 496 3161
rect -496 3121 496 3127
rect -496 3053 496 3059
rect -496 3019 -484 3053
rect 484 3019 496 3053
rect -496 3013 496 3019
rect -552 2960 -506 2972
rect -552 1984 -546 2960
rect -512 1984 -506 2960
rect -552 1972 -506 1984
rect 506 2960 552 2972
rect 506 1984 512 2960
rect 546 1984 552 2960
rect 506 1972 552 1984
rect -496 1925 496 1931
rect -496 1891 -484 1925
rect 484 1891 496 1925
rect -496 1885 496 1891
rect -496 1817 496 1823
rect -496 1783 -484 1817
rect 484 1783 496 1817
rect -496 1777 496 1783
rect -552 1724 -506 1736
rect -552 748 -546 1724
rect -512 748 -506 1724
rect -552 736 -506 748
rect 506 1724 552 1736
rect 506 748 512 1724
rect 546 748 552 1724
rect 506 736 552 748
rect -496 689 496 695
rect -496 655 -484 689
rect 484 655 496 689
rect -496 649 496 655
rect -496 581 496 587
rect -496 547 -484 581
rect 484 547 496 581
rect -496 541 496 547
rect -552 488 -506 500
rect -552 -488 -546 488
rect -512 -488 -506 488
rect -552 -500 -506 -488
rect 506 488 552 500
rect 506 -488 512 488
rect 546 -488 552 488
rect 506 -500 552 -488
rect -496 -547 496 -541
rect -496 -581 -484 -547
rect 484 -581 496 -547
rect -496 -587 496 -581
rect -496 -655 496 -649
rect -496 -689 -484 -655
rect 484 -689 496 -655
rect -496 -695 496 -689
rect -552 -748 -506 -736
rect -552 -1724 -546 -748
rect -512 -1724 -506 -748
rect -552 -1736 -506 -1724
rect 506 -748 552 -736
rect 506 -1724 512 -748
rect 546 -1724 552 -748
rect 506 -1736 552 -1724
rect -496 -1783 496 -1777
rect -496 -1817 -484 -1783
rect 484 -1817 496 -1783
rect -496 -1823 496 -1817
rect -496 -1891 496 -1885
rect -496 -1925 -484 -1891
rect 484 -1925 496 -1891
rect -496 -1931 496 -1925
rect -552 -1984 -506 -1972
rect -552 -2960 -546 -1984
rect -512 -2960 -506 -1984
rect -552 -2972 -506 -2960
rect 506 -1984 552 -1972
rect 506 -2960 512 -1984
rect 546 -2960 552 -1984
rect 506 -2972 552 -2960
rect -496 -3019 496 -3013
rect -496 -3053 -484 -3019
rect 484 -3053 496 -3019
rect -496 -3059 496 -3053
rect -496 -3127 496 -3121
rect -496 -3161 -484 -3127
rect 484 -3161 496 -3127
rect -496 -3167 496 -3161
rect -552 -3220 -506 -3208
rect -552 -4196 -546 -3220
rect -512 -4196 -506 -3220
rect -552 -4208 -506 -4196
rect 506 -3220 552 -3208
rect 506 -4196 512 -3220
rect 546 -4196 552 -3220
rect 506 -4208 552 -4196
rect -496 -4255 496 -4249
rect -496 -4289 -484 -4255
rect 484 -4289 496 -4255
rect -496 -4295 496 -4289
rect -496 -4363 496 -4357
rect -496 -4397 -484 -4363
rect 484 -4397 496 -4363
rect -496 -4403 496 -4397
rect -552 -4456 -506 -4444
rect -552 -5432 -546 -4456
rect -512 -5432 -506 -4456
rect -552 -5444 -506 -5432
rect 506 -4456 552 -4444
rect 506 -5432 512 -4456
rect 546 -5432 552 -4456
rect 506 -5444 552 -5432
rect -496 -5491 496 -5485
rect -496 -5525 -484 -5491
rect 484 -5525 496 -5491
rect -496 -5531 496 -5525
rect -496 -5599 496 -5593
rect -496 -5633 -484 -5599
rect 484 -5633 496 -5599
rect -496 -5639 496 -5633
rect -552 -5692 -506 -5680
rect -552 -6668 -546 -5692
rect -512 -6668 -506 -5692
rect -552 -6680 -506 -6668
rect 506 -5692 552 -5680
rect 506 -6668 512 -5692
rect 546 -6668 552 -5692
rect 506 -6680 552 -6668
rect -496 -6727 496 -6721
rect -496 -6761 -484 -6727
rect 484 -6761 496 -6727
rect -496 -6767 496 -6761
rect -496 -6835 496 -6829
rect -496 -6869 -484 -6835
rect 484 -6869 496 -6835
rect -496 -6875 496 -6869
rect -552 -6928 -506 -6916
rect -552 -7904 -546 -6928
rect -512 -7904 -506 -6928
rect -552 -7916 -506 -7904
rect 506 -6928 552 -6916
rect 506 -7904 512 -6928
rect 546 -7904 552 -6928
rect 506 -7916 552 -7904
rect -496 -7963 496 -7957
rect -496 -7997 -484 -7963
rect 484 -7997 496 -7963
rect -496 -8003 496 -7997
rect -496 -8071 496 -8065
rect -496 -8105 -484 -8071
rect 484 -8105 496 -8071
rect -496 -8111 496 -8105
rect -552 -8164 -506 -8152
rect -552 -9140 -546 -8164
rect -512 -9140 -506 -8164
rect -552 -9152 -506 -9140
rect 506 -8164 552 -8152
rect 506 -9140 512 -8164
rect 546 -9140 552 -8164
rect 506 -9152 552 -9140
rect -496 -9199 496 -9193
rect -496 -9233 -484 -9199
rect 484 -9233 496 -9199
rect -496 -9239 496 -9233
<< properties >>
string FIXED_BBOX -643 -9318 643 9318
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 5.0 l 5.0 m 15 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
