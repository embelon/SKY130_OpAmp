magic
tech sky130A
magscale 1 2
timestamp 1695666882
<< nmos >>
rect -100 1045 100 1295
rect -100 577 100 827
rect -100 109 100 359
rect -100 -359 100 -109
rect -100 -827 100 -577
rect -100 -1295 100 -1045
<< ndiff >>
rect -158 1283 -100 1295
rect -158 1057 -146 1283
rect -112 1057 -100 1283
rect -158 1045 -100 1057
rect 100 1283 158 1295
rect 100 1057 112 1283
rect 146 1057 158 1283
rect 100 1045 158 1057
rect -158 815 -100 827
rect -158 589 -146 815
rect -112 589 -100 815
rect -158 577 -100 589
rect 100 815 158 827
rect 100 589 112 815
rect 146 589 158 815
rect 100 577 158 589
rect -158 347 -100 359
rect -158 121 -146 347
rect -112 121 -100 347
rect -158 109 -100 121
rect 100 347 158 359
rect 100 121 112 347
rect 146 121 158 347
rect 100 109 158 121
rect -158 -121 -100 -109
rect -158 -347 -146 -121
rect -112 -347 -100 -121
rect -158 -359 -100 -347
rect 100 -121 158 -109
rect 100 -347 112 -121
rect 146 -347 158 -121
rect 100 -359 158 -347
rect -158 -589 -100 -577
rect -158 -815 -146 -589
rect -112 -815 -100 -589
rect -158 -827 -100 -815
rect 100 -589 158 -577
rect 100 -815 112 -589
rect 146 -815 158 -589
rect 100 -827 158 -815
rect -158 -1057 -100 -1045
rect -158 -1283 -146 -1057
rect -112 -1283 -100 -1057
rect -158 -1295 -100 -1283
rect 100 -1057 158 -1045
rect 100 -1283 112 -1057
rect 146 -1283 158 -1057
rect 100 -1295 158 -1283
<< ndiffc >>
rect -146 1057 -112 1283
rect 112 1057 146 1283
rect -146 589 -112 815
rect 112 589 146 815
rect -146 121 -112 347
rect 112 121 146 347
rect -146 -347 -112 -121
rect 112 -347 146 -121
rect -146 -815 -112 -589
rect 112 -815 146 -589
rect -146 -1283 -112 -1057
rect 112 -1283 146 -1057
<< poly >>
rect -100 1367 100 1383
rect -100 1333 -84 1367
rect 84 1333 100 1367
rect -100 1295 100 1333
rect -100 1007 100 1045
rect -100 973 -84 1007
rect 84 973 100 1007
rect -100 957 100 973
rect -100 899 100 915
rect -100 865 -84 899
rect 84 865 100 899
rect -100 827 100 865
rect -100 539 100 577
rect -100 505 -84 539
rect 84 505 100 539
rect -100 489 100 505
rect -100 431 100 447
rect -100 397 -84 431
rect 84 397 100 431
rect -100 359 100 397
rect -100 71 100 109
rect -100 37 -84 71
rect 84 37 100 71
rect -100 21 100 37
rect -100 -37 100 -21
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -100 -109 100 -71
rect -100 -397 100 -359
rect -100 -431 -84 -397
rect 84 -431 100 -397
rect -100 -447 100 -431
rect -100 -505 100 -489
rect -100 -539 -84 -505
rect 84 -539 100 -505
rect -100 -577 100 -539
rect -100 -865 100 -827
rect -100 -899 -84 -865
rect 84 -899 100 -865
rect -100 -915 100 -899
rect -100 -973 100 -957
rect -100 -1007 -84 -973
rect 84 -1007 100 -973
rect -100 -1045 100 -1007
rect -100 -1333 100 -1295
rect -100 -1367 -84 -1333
rect 84 -1367 100 -1333
rect -100 -1383 100 -1367
<< polycont >>
rect -84 1333 84 1367
rect -84 973 84 1007
rect -84 865 84 899
rect -84 505 84 539
rect -84 397 84 431
rect -84 37 84 71
rect -84 -71 84 -37
rect -84 -431 84 -397
rect -84 -539 84 -505
rect -84 -899 84 -865
rect -84 -1007 84 -973
rect -84 -1367 84 -1333
<< locali >>
rect -100 1333 -84 1367
rect 84 1333 100 1367
rect -146 1283 -112 1299
rect -146 1041 -112 1057
rect 112 1283 146 1299
rect 112 1041 146 1057
rect -100 973 -84 1007
rect 84 973 100 1007
rect -100 865 -84 899
rect 84 865 100 899
rect -146 815 -112 831
rect -146 573 -112 589
rect 112 815 146 831
rect 112 573 146 589
rect -100 505 -84 539
rect 84 505 100 539
rect -100 397 -84 431
rect 84 397 100 431
rect -146 347 -112 363
rect -146 105 -112 121
rect 112 347 146 363
rect 112 105 146 121
rect -100 37 -84 71
rect 84 37 100 71
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -146 -121 -112 -105
rect -146 -363 -112 -347
rect 112 -121 146 -105
rect 112 -363 146 -347
rect -100 -431 -84 -397
rect 84 -431 100 -397
rect -100 -539 -84 -505
rect 84 -539 100 -505
rect -146 -589 -112 -573
rect -146 -831 -112 -815
rect 112 -589 146 -573
rect 112 -831 146 -815
rect -100 -899 -84 -865
rect 84 -899 100 -865
rect -100 -1007 -84 -973
rect 84 -1007 100 -973
rect -146 -1057 -112 -1041
rect -146 -1299 -112 -1283
rect 112 -1057 146 -1041
rect 112 -1299 146 -1283
rect -100 -1367 -84 -1333
rect 84 -1367 100 -1333
<< viali >>
rect -84 1333 84 1367
rect -146 1057 -112 1283
rect 112 1057 146 1283
rect -84 973 84 1007
rect -84 865 84 899
rect -146 589 -112 815
rect 112 589 146 815
rect -84 505 84 539
rect -84 397 84 431
rect -146 121 -112 347
rect 112 121 146 347
rect -84 37 84 71
rect -84 -71 84 -37
rect -146 -347 -112 -121
rect 112 -347 146 -121
rect -84 -431 84 -397
rect -84 -539 84 -505
rect -146 -815 -112 -589
rect 112 -815 146 -589
rect -84 -899 84 -865
rect -84 -1007 84 -973
rect -146 -1283 -112 -1057
rect 112 -1283 146 -1057
rect -84 -1367 84 -1333
<< metal1 >>
rect -96 1367 96 1373
rect -96 1333 -84 1367
rect 84 1333 96 1367
rect -96 1327 96 1333
rect -152 1283 -106 1295
rect -152 1057 -146 1283
rect -112 1057 -106 1283
rect -152 1045 -106 1057
rect 106 1283 152 1295
rect 106 1057 112 1283
rect 146 1057 152 1283
rect 106 1045 152 1057
rect -96 1007 96 1013
rect -96 973 -84 1007
rect 84 973 96 1007
rect -96 967 96 973
rect -96 899 96 905
rect -96 865 -84 899
rect 84 865 96 899
rect -96 859 96 865
rect -152 815 -106 827
rect -152 589 -146 815
rect -112 589 -106 815
rect -152 577 -106 589
rect 106 815 152 827
rect 106 589 112 815
rect 146 589 152 815
rect 106 577 152 589
rect -96 539 96 545
rect -96 505 -84 539
rect 84 505 96 539
rect -96 499 96 505
rect -96 431 96 437
rect -96 397 -84 431
rect 84 397 96 431
rect -96 391 96 397
rect -152 347 -106 359
rect -152 121 -146 347
rect -112 121 -106 347
rect -152 109 -106 121
rect 106 347 152 359
rect 106 121 112 347
rect 146 121 152 347
rect 106 109 152 121
rect -96 71 96 77
rect -96 37 -84 71
rect 84 37 96 71
rect -96 31 96 37
rect -96 -37 96 -31
rect -96 -71 -84 -37
rect 84 -71 96 -37
rect -96 -77 96 -71
rect -152 -121 -106 -109
rect -152 -347 -146 -121
rect -112 -347 -106 -121
rect -152 -359 -106 -347
rect 106 -121 152 -109
rect 106 -347 112 -121
rect 146 -347 152 -121
rect 106 -359 152 -347
rect -96 -397 96 -391
rect -96 -431 -84 -397
rect 84 -431 96 -397
rect -96 -437 96 -431
rect -96 -505 96 -499
rect -96 -539 -84 -505
rect 84 -539 96 -505
rect -96 -545 96 -539
rect -152 -589 -106 -577
rect -152 -815 -146 -589
rect -112 -815 -106 -589
rect -152 -827 -106 -815
rect 106 -589 152 -577
rect 106 -815 112 -589
rect 146 -815 152 -589
rect 106 -827 152 -815
rect -96 -865 96 -859
rect -96 -899 -84 -865
rect 84 -899 96 -865
rect -96 -905 96 -899
rect -96 -973 96 -967
rect -96 -1007 -84 -973
rect 84 -1007 96 -973
rect -96 -1013 96 -1007
rect -152 -1057 -106 -1045
rect -152 -1283 -146 -1057
rect -112 -1283 -106 -1057
rect -152 -1295 -106 -1283
rect 106 -1057 152 -1045
rect 106 -1283 112 -1057
rect 146 -1283 152 -1057
rect 106 -1295 152 -1283
rect -96 -1333 96 -1327
rect -96 -1367 -84 -1333
rect 84 -1367 96 -1333
rect -96 -1373 96 -1367
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.25 l 1 m 6 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
