** sch_path: ../opamp_cascode_dc_max_gain.sch
**.subckt opamp_cascode_dc_max_gain
Vcm net1 GND 0.9
.save i(vcm)
C1 out GND 1p m=1
Vdiff Vdiff GND 0
.save i(vdiff)
Ib IBIAS GND 45u
B1 Vp net1 v=v(Vdiff)
B2 net1 Vn v=v(Vdiff)
x1 Vp Vn VCC GND out VB_A VB_B IBIAS opamp_cascode
**** begin user architecture code


Vsupply VCC GND 1.8
VbiasA VB_A GND 0.2
VbiasB VB_B GND 1.1
.include ../opamp_cascode.spice
.control
  save all
  dc Vdiff -0.01 0.01 0.000001
  let dVout = deriv(v(out))
  plot dVout vs Vdiff retraceplot
  meas dc maxGain max dVout
  set hcopydevtype = svg
  hardcopy dc_max_gain.svg dVout vs Vdiff
.endc



.param mc_mm_switch=1
.param mc_pr_switch=0
.include ~/.volare/sky130A/libs.tech/ngspice/corners/tt.spice
.include ~/.volare/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include ~/.volare/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include ~/.volare/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice

**** end user architecture code
**.ends
.GLOBAL GND
.end
