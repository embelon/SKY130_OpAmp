magic
tech sky130A
magscale 1 2
timestamp 1695661682
<< nwell >>
rect -496 -1955 496 1955
<< pmos >>
rect -300 736 300 1736
rect -300 -500 300 500
rect -300 -1736 300 -736
<< pdiff >>
rect -358 1724 -300 1736
rect -358 748 -346 1724
rect -312 748 -300 1724
rect -358 736 -300 748
rect 300 1724 358 1736
rect 300 748 312 1724
rect 346 748 358 1724
rect 300 736 358 748
rect -358 488 -300 500
rect -358 -488 -346 488
rect -312 -488 -300 488
rect -358 -500 -300 -488
rect 300 488 358 500
rect 300 -488 312 488
rect 346 -488 358 488
rect 300 -500 358 -488
rect -358 -748 -300 -736
rect -358 -1724 -346 -748
rect -312 -1724 -300 -748
rect -358 -1736 -300 -1724
rect 300 -748 358 -736
rect 300 -1724 312 -748
rect 346 -1724 358 -748
rect 300 -1736 358 -1724
<< pdiffc >>
rect -346 748 -312 1724
rect 312 748 346 1724
rect -346 -488 -312 488
rect 312 -488 346 488
rect -346 -1724 -312 -748
rect 312 -1724 346 -748
<< nsubdiff >>
rect -460 1885 -364 1919
rect 364 1885 460 1919
rect -460 1823 -426 1885
rect 426 1823 460 1885
rect -460 -1885 -426 -1823
rect 426 -1885 460 -1823
rect -460 -1919 -364 -1885
rect 364 -1919 460 -1885
<< nsubdiffcont >>
rect -364 1885 364 1919
rect -460 -1823 -426 1823
rect 426 -1823 460 1823
rect -364 -1919 364 -1885
<< poly >>
rect -300 1817 300 1833
rect -300 1783 -284 1817
rect 284 1783 300 1817
rect -300 1736 300 1783
rect -300 689 300 736
rect -300 655 -284 689
rect 284 655 300 689
rect -300 639 300 655
rect -300 581 300 597
rect -300 547 -284 581
rect 284 547 300 581
rect -300 500 300 547
rect -300 -547 300 -500
rect -300 -581 -284 -547
rect 284 -581 300 -547
rect -300 -597 300 -581
rect -300 -655 300 -639
rect -300 -689 -284 -655
rect 284 -689 300 -655
rect -300 -736 300 -689
rect -300 -1783 300 -1736
rect -300 -1817 -284 -1783
rect 284 -1817 300 -1783
rect -300 -1833 300 -1817
<< polycont >>
rect -284 1783 284 1817
rect -284 655 284 689
rect -284 547 284 581
rect -284 -581 284 -547
rect -284 -689 284 -655
rect -284 -1817 284 -1783
<< locali >>
rect -460 1885 -364 1919
rect 364 1885 460 1919
rect -460 1823 -426 1885
rect 426 1823 460 1885
rect -300 1783 -284 1817
rect 284 1783 300 1817
rect -346 1724 -312 1740
rect -346 732 -312 748
rect 312 1724 346 1740
rect 312 732 346 748
rect -300 655 -284 689
rect 284 655 300 689
rect -300 547 -284 581
rect 284 547 300 581
rect -346 488 -312 504
rect -346 -504 -312 -488
rect 312 488 346 504
rect 312 -504 346 -488
rect -300 -581 -284 -547
rect 284 -581 300 -547
rect -300 -689 -284 -655
rect 284 -689 300 -655
rect -346 -748 -312 -732
rect -346 -1740 -312 -1724
rect 312 -748 346 -732
rect 312 -1740 346 -1724
rect -300 -1817 -284 -1783
rect 284 -1817 300 -1783
rect -460 -1885 -426 -1823
rect 426 -1885 460 -1823
rect -460 -1919 -364 -1885
rect 364 -1919 460 -1885
<< viali >>
rect -284 1783 284 1817
rect -346 748 -312 1724
rect 312 748 346 1724
rect -284 655 284 689
rect -284 547 284 581
rect -346 -488 -312 488
rect 312 -488 346 488
rect -284 -581 284 -547
rect -284 -689 284 -655
rect -346 -1724 -312 -748
rect 312 -1724 346 -748
rect -284 -1817 284 -1783
<< metal1 >>
rect -296 1817 296 1823
rect -296 1783 -284 1817
rect 284 1783 296 1817
rect -296 1777 296 1783
rect -352 1724 -306 1736
rect -352 748 -346 1724
rect -312 748 -306 1724
rect -352 736 -306 748
rect 306 1724 352 1736
rect 306 748 312 1724
rect 346 748 352 1724
rect 306 736 352 748
rect -296 689 296 695
rect -296 655 -284 689
rect 284 655 296 689
rect -296 649 296 655
rect -296 581 296 587
rect -296 547 -284 581
rect 284 547 296 581
rect -296 541 296 547
rect -352 488 -306 500
rect -352 -488 -346 488
rect -312 -488 -306 488
rect -352 -500 -306 -488
rect 306 488 352 500
rect 306 -488 312 488
rect 346 -488 352 488
rect 306 -500 352 -488
rect -296 -547 296 -541
rect -296 -581 -284 -547
rect 284 -581 296 -547
rect -296 -587 296 -581
rect -296 -655 296 -649
rect -296 -689 -284 -655
rect 284 -689 296 -655
rect -296 -695 296 -689
rect -352 -748 -306 -736
rect -352 -1724 -346 -748
rect -312 -1724 -306 -748
rect -352 -1736 -306 -1724
rect 306 -748 352 -736
rect 306 -1724 312 -748
rect 346 -1724 352 -748
rect 306 -1736 352 -1724
rect -296 -1783 296 -1777
rect -296 -1817 -284 -1783
rect 284 -1817 296 -1783
rect -296 -1823 296 -1817
<< properties >>
string FIXED_BBOX -443 -1902 443 1902
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 5.0 l 3.0 m 3 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
