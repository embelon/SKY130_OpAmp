** sch_path: /home/zwierzak/projects/SKY130_OpAmp/06_ParasiticsSim/opamp_cascode_ac_psrr.sch
**.subckt opamp_cascode_ac_psrr
C1 out GND 1p m=1
x1 VCC GND VB_B Vcm Vn out IBIAS VB_A opamp_cascode
I0 IBIAS GND 45u
R1 out Vn 1k m=1
V1 Vcm GND 0.9
.save i(v1)
**** begin user architecture code


Vsupply VCC GND 1.8
VbiasA VB_A GND 0.2
VbiasB VB_B GND 1.1
.include ../opamp_cascode.spice
.control
  alter Vsupply AC = 1
  save all
  ac dec 10 1 1G
  let invVn = 1/(v(Vcm)-v(Vn))
  plot db(invVn)
  meas ac PSR_1k FIND vdb(invVn) AT=1k
  meas ac PSR_1M FIND vdb(invVn) AT=1Meg
  echo PSRR_1k = $&PSR_1k dB
  echo PSRR_1M = $&PSR_1M dB
.endc



.param mc_mm_switch=0
.param mc_pr_switch=0
.include ~/.volare/sky130A/libs.tech/ngspice/corners/tt.spice
.include ~/.volare/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include ~/.volare/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include ~/.volare/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice

**** end user architecture code
**.ends
.GLOBAL GND
.end
