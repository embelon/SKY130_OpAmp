VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO opamp_cascode
  CLASS BLOCK ;
  FOREIGN opamp_cascode ;
  ORIGIN -181.000 -70.000 ;
  SIZE 349.000 BY 655.050 ;
  PIN IN_P
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 64.799995 ;
    PORT
      LAYER met3 ;
        RECT 181.000 72.000 185.000 74.000 ;
    END
  END IN_P
  PIN IN_M
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 27.000000 ;
    PORT
      LAYER met3 ;
        RECT 181.000 76.000 185.000 78.000 ;
    END
  END IN_M
  PIN VCC
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 190.000 248.000 200.000 725.000 ;
    END
  END VCC
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 267.000 684.000 277.000 725.000 ;
    END
  END VSS
  PIN OUT
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 87.000000 ;
    PORT
      LAYER met3 ;
        RECT 181.000 452.000 185.000 454.000 ;
    END
  END OUT
  PIN VB_A
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2550.000000 ;
    PORT
      LAYER met3 ;
        RECT 181.000 437.000 185.000 439.000 ;
    END
  END VB_A
  PIN VB_B
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2550.000000 ;
    PORT
      LAYER met3 ;
        RECT 181.000 564.000 185.000 566.000 ;
    END
  END VB_B
  PIN IB
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 450.000000 ;
    ANTENNADIFFAREA 5.800000 ;
    PORT
      LAYER met3 ;
        RECT 181.000 271.000 185.000 273.000 ;
    END
  END IB
  OBS
      LAYER li1 ;
        RECT 218.060 79.095 523.700 719.400 ;
      LAYER met1 ;
        RECT 205.950 74.500 524.500 725.000 ;
      LAYER met2 ;
        RECT 186.000 71.950 524.000 725.050 ;
      LAYER met3 ;
        RECT 185.000 566.400 277.000 725.000 ;
        RECT 185.400 563.600 277.000 566.400 ;
        RECT 185.000 454.400 277.000 563.600 ;
        RECT 185.400 451.600 277.000 454.400 ;
        RECT 185.000 439.400 277.000 451.600 ;
        RECT 185.400 436.600 277.000 439.400 ;
        RECT 185.000 273.400 277.000 436.600 ;
        RECT 185.400 270.600 277.000 273.400 ;
        RECT 185.000 78.400 277.000 270.600 ;
        RECT 185.400 75.600 277.000 78.400 ;
        RECT 185.000 74.400 277.000 75.600 ;
        RECT 185.400 71.975 277.000 74.400 ;
      LAYER met4 ;
        RECT 200.400 683.600 266.600 725.000 ;
        RECT 200.400 247.600 277.000 683.600 ;
        RECT 190.000 246.000 277.000 247.600 ;
  END
END opamp_cascode
END LIBRARY

