magic
tech sky130A
magscale 1 2
timestamp 1695661682
<< pwell >>
rect -321 -1355 321 1355
<< nmos >>
rect -125 945 125 1145
rect -125 527 125 727
rect -125 109 125 309
rect -125 -309 125 -109
rect -125 -727 125 -527
rect -125 -1145 125 -945
<< ndiff >>
rect -183 1133 -125 1145
rect -183 957 -171 1133
rect -137 957 -125 1133
rect -183 945 -125 957
rect 125 1133 183 1145
rect 125 957 137 1133
rect 171 957 183 1133
rect 125 945 183 957
rect -183 715 -125 727
rect -183 539 -171 715
rect -137 539 -125 715
rect -183 527 -125 539
rect 125 715 183 727
rect 125 539 137 715
rect 171 539 183 715
rect 125 527 183 539
rect -183 297 -125 309
rect -183 121 -171 297
rect -137 121 -125 297
rect -183 109 -125 121
rect 125 297 183 309
rect 125 121 137 297
rect 171 121 183 297
rect 125 109 183 121
rect -183 -121 -125 -109
rect -183 -297 -171 -121
rect -137 -297 -125 -121
rect -183 -309 -125 -297
rect 125 -121 183 -109
rect 125 -297 137 -121
rect 171 -297 183 -121
rect 125 -309 183 -297
rect -183 -539 -125 -527
rect -183 -715 -171 -539
rect -137 -715 -125 -539
rect -183 -727 -125 -715
rect 125 -539 183 -527
rect 125 -715 137 -539
rect 171 -715 183 -539
rect 125 -727 183 -715
rect -183 -957 -125 -945
rect -183 -1133 -171 -957
rect -137 -1133 -125 -957
rect -183 -1145 -125 -1133
rect 125 -957 183 -945
rect 125 -1133 137 -957
rect 171 -1133 183 -957
rect 125 -1145 183 -1133
<< ndiffc >>
rect -171 957 -137 1133
rect 137 957 171 1133
rect -171 539 -137 715
rect 137 539 171 715
rect -171 121 -137 297
rect 137 121 171 297
rect -171 -297 -137 -121
rect 137 -297 171 -121
rect -171 -715 -137 -539
rect 137 -715 171 -539
rect -171 -1133 -137 -957
rect 137 -1133 171 -957
<< psubdiff >>
rect -285 1285 -189 1319
rect 189 1285 285 1319
rect -285 1223 -251 1285
rect 251 1223 285 1285
rect -285 -1285 -251 -1223
rect 251 -1285 285 -1223
rect -285 -1319 -189 -1285
rect 189 -1319 285 -1285
<< psubdiffcont >>
rect -189 1285 189 1319
rect -285 -1223 -251 1223
rect 251 -1223 285 1223
rect -189 -1319 189 -1285
<< poly >>
rect -125 1217 125 1233
rect -125 1183 -109 1217
rect 109 1183 125 1217
rect -125 1145 125 1183
rect -125 907 125 945
rect -125 873 -109 907
rect 109 873 125 907
rect -125 857 125 873
rect -125 799 125 815
rect -125 765 -109 799
rect 109 765 125 799
rect -125 727 125 765
rect -125 489 125 527
rect -125 455 -109 489
rect 109 455 125 489
rect -125 439 125 455
rect -125 381 125 397
rect -125 347 -109 381
rect 109 347 125 381
rect -125 309 125 347
rect -125 71 125 109
rect -125 37 -109 71
rect 109 37 125 71
rect -125 21 125 37
rect -125 -37 125 -21
rect -125 -71 -109 -37
rect 109 -71 125 -37
rect -125 -109 125 -71
rect -125 -347 125 -309
rect -125 -381 -109 -347
rect 109 -381 125 -347
rect -125 -397 125 -381
rect -125 -455 125 -439
rect -125 -489 -109 -455
rect 109 -489 125 -455
rect -125 -527 125 -489
rect -125 -765 125 -727
rect -125 -799 -109 -765
rect 109 -799 125 -765
rect -125 -815 125 -799
rect -125 -873 125 -857
rect -125 -907 -109 -873
rect 109 -907 125 -873
rect -125 -945 125 -907
rect -125 -1183 125 -1145
rect -125 -1217 -109 -1183
rect 109 -1217 125 -1183
rect -125 -1233 125 -1217
<< polycont >>
rect -109 1183 109 1217
rect -109 873 109 907
rect -109 765 109 799
rect -109 455 109 489
rect -109 347 109 381
rect -109 37 109 71
rect -109 -71 109 -37
rect -109 -381 109 -347
rect -109 -489 109 -455
rect -109 -799 109 -765
rect -109 -907 109 -873
rect -109 -1217 109 -1183
<< locali >>
rect -285 1285 -189 1319
rect 189 1285 285 1319
rect -285 1223 -251 1285
rect 251 1223 285 1285
rect -125 1183 -109 1217
rect 109 1183 125 1217
rect -171 1133 -137 1149
rect -171 941 -137 957
rect 137 1133 171 1149
rect 137 941 171 957
rect -125 873 -109 907
rect 109 873 125 907
rect -125 765 -109 799
rect 109 765 125 799
rect -171 715 -137 731
rect -171 523 -137 539
rect 137 715 171 731
rect 137 523 171 539
rect -125 455 -109 489
rect 109 455 125 489
rect -125 347 -109 381
rect 109 347 125 381
rect -171 297 -137 313
rect -171 105 -137 121
rect 137 297 171 313
rect 137 105 171 121
rect -125 37 -109 71
rect 109 37 125 71
rect -125 -71 -109 -37
rect 109 -71 125 -37
rect -171 -121 -137 -105
rect -171 -313 -137 -297
rect 137 -121 171 -105
rect 137 -313 171 -297
rect -125 -381 -109 -347
rect 109 -381 125 -347
rect -125 -489 -109 -455
rect 109 -489 125 -455
rect -171 -539 -137 -523
rect -171 -731 -137 -715
rect 137 -539 171 -523
rect 137 -731 171 -715
rect -125 -799 -109 -765
rect 109 -799 125 -765
rect -125 -907 -109 -873
rect 109 -907 125 -873
rect -171 -957 -137 -941
rect -171 -1149 -137 -1133
rect 137 -957 171 -941
rect 137 -1149 171 -1133
rect -125 -1217 -109 -1183
rect 109 -1217 125 -1183
rect -285 -1285 -251 -1223
rect 251 -1285 285 -1223
rect -285 -1319 -189 -1285
rect 189 -1319 285 -1285
<< viali >>
rect -109 1183 109 1217
rect -171 957 -137 1133
rect 137 957 171 1133
rect -109 873 109 907
rect -109 765 109 799
rect -171 539 -137 715
rect 137 539 171 715
rect -109 455 109 489
rect -109 347 109 381
rect -171 121 -137 297
rect 137 121 171 297
rect -109 37 109 71
rect -109 -71 109 -37
rect -171 -297 -137 -121
rect 137 -297 171 -121
rect -109 -381 109 -347
rect -109 -489 109 -455
rect -171 -715 -137 -539
rect 137 -715 171 -539
rect -109 -799 109 -765
rect -109 -907 109 -873
rect -171 -1133 -137 -957
rect 137 -1133 171 -957
rect -109 -1217 109 -1183
<< metal1 >>
rect -121 1217 121 1223
rect -121 1183 -109 1217
rect 109 1183 121 1217
rect -121 1177 121 1183
rect -177 1133 -131 1145
rect -177 957 -171 1133
rect -137 957 -131 1133
rect -177 945 -131 957
rect 131 1133 177 1145
rect 131 957 137 1133
rect 171 957 177 1133
rect 131 945 177 957
rect -121 907 121 913
rect -121 873 -109 907
rect 109 873 121 907
rect -121 867 121 873
rect -121 799 121 805
rect -121 765 -109 799
rect 109 765 121 799
rect -121 759 121 765
rect -177 715 -131 727
rect -177 539 -171 715
rect -137 539 -131 715
rect -177 527 -131 539
rect 131 715 177 727
rect 131 539 137 715
rect 171 539 177 715
rect 131 527 177 539
rect -121 489 121 495
rect -121 455 -109 489
rect 109 455 121 489
rect -121 449 121 455
rect -121 381 121 387
rect -121 347 -109 381
rect 109 347 121 381
rect -121 341 121 347
rect -177 297 -131 309
rect -177 121 -171 297
rect -137 121 -131 297
rect -177 109 -131 121
rect 131 297 177 309
rect 131 121 137 297
rect 171 121 177 297
rect 131 109 177 121
rect -121 71 121 77
rect -121 37 -109 71
rect 109 37 121 71
rect -121 31 121 37
rect -121 -37 121 -31
rect -121 -71 -109 -37
rect 109 -71 121 -37
rect -121 -77 121 -71
rect -177 -121 -131 -109
rect -177 -297 -171 -121
rect -137 -297 -131 -121
rect -177 -309 -131 -297
rect 131 -121 177 -109
rect 131 -297 137 -121
rect 171 -297 177 -121
rect 131 -309 177 -297
rect -121 -347 121 -341
rect -121 -381 -109 -347
rect 109 -381 121 -347
rect -121 -387 121 -381
rect -121 -455 121 -449
rect -121 -489 -109 -455
rect 109 -489 121 -455
rect -121 -495 121 -489
rect -177 -539 -131 -527
rect -177 -715 -171 -539
rect -137 -715 -131 -539
rect -177 -727 -131 -715
rect 131 -539 177 -527
rect 131 -715 137 -539
rect 171 -715 177 -539
rect 131 -727 177 -715
rect -121 -765 121 -759
rect -121 -799 -109 -765
rect 109 -799 121 -765
rect -121 -805 121 -799
rect -121 -873 121 -867
rect -121 -907 -109 -873
rect 109 -907 121 -873
rect -121 -913 121 -907
rect -177 -957 -131 -945
rect -177 -1133 -171 -957
rect -137 -1133 -131 -957
rect -177 -1145 -131 -1133
rect 131 -957 177 -945
rect 131 -1133 137 -957
rect 171 -1133 177 -957
rect 131 -1145 177 -1133
rect -121 -1183 121 -1177
rect -121 -1217 -109 -1183
rect 109 -1217 121 -1183
rect -121 -1223 121 -1217
<< properties >>
string FIXED_BBOX -268 -1302 268 1302
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.0 l 1.25 m 6 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
