magic
tech sky130A
timestamp 1695666081
<< nmos >>
rect -250 4013 250 4513
rect -250 3404 250 3904
rect -250 2795 250 3295
rect -250 2186 250 2686
rect -250 1577 250 2077
rect -250 968 250 1468
rect -250 359 250 859
rect -250 -250 250 250
rect -250 -859 250 -359
rect -250 -1468 250 -968
rect -250 -2077 250 -1577
rect -250 -2686 250 -2186
rect -250 -3295 250 -2795
rect -250 -3904 250 -3404
rect -250 -4513 250 -4013
<< ndiff >>
rect -279 4507 -250 4513
rect -279 4019 -273 4507
rect -256 4019 -250 4507
rect -279 4013 -250 4019
rect 250 4507 279 4513
rect 250 4019 256 4507
rect 273 4019 279 4507
rect 250 4013 279 4019
rect -279 3898 -250 3904
rect -279 3410 -273 3898
rect -256 3410 -250 3898
rect -279 3404 -250 3410
rect 250 3898 279 3904
rect 250 3410 256 3898
rect 273 3410 279 3898
rect 250 3404 279 3410
rect -279 3289 -250 3295
rect -279 2801 -273 3289
rect -256 2801 -250 3289
rect -279 2795 -250 2801
rect 250 3289 279 3295
rect 250 2801 256 3289
rect 273 2801 279 3289
rect 250 2795 279 2801
rect -279 2680 -250 2686
rect -279 2192 -273 2680
rect -256 2192 -250 2680
rect -279 2186 -250 2192
rect 250 2680 279 2686
rect 250 2192 256 2680
rect 273 2192 279 2680
rect 250 2186 279 2192
rect -279 2071 -250 2077
rect -279 1583 -273 2071
rect -256 1583 -250 2071
rect -279 1577 -250 1583
rect 250 2071 279 2077
rect 250 1583 256 2071
rect 273 1583 279 2071
rect 250 1577 279 1583
rect -279 1462 -250 1468
rect -279 974 -273 1462
rect -256 974 -250 1462
rect -279 968 -250 974
rect 250 1462 279 1468
rect 250 974 256 1462
rect 273 974 279 1462
rect 250 968 279 974
rect -279 853 -250 859
rect -279 365 -273 853
rect -256 365 -250 853
rect -279 359 -250 365
rect 250 853 279 859
rect 250 365 256 853
rect 273 365 279 853
rect 250 359 279 365
rect -279 244 -250 250
rect -279 -244 -273 244
rect -256 -244 -250 244
rect -279 -250 -250 -244
rect 250 244 279 250
rect 250 -244 256 244
rect 273 -244 279 244
rect 250 -250 279 -244
rect -279 -365 -250 -359
rect -279 -853 -273 -365
rect -256 -853 -250 -365
rect -279 -859 -250 -853
rect 250 -365 279 -359
rect 250 -853 256 -365
rect 273 -853 279 -365
rect 250 -859 279 -853
rect -279 -974 -250 -968
rect -279 -1462 -273 -974
rect -256 -1462 -250 -974
rect -279 -1468 -250 -1462
rect 250 -974 279 -968
rect 250 -1462 256 -974
rect 273 -1462 279 -974
rect 250 -1468 279 -1462
rect -279 -1583 -250 -1577
rect -279 -2071 -273 -1583
rect -256 -2071 -250 -1583
rect -279 -2077 -250 -2071
rect 250 -1583 279 -1577
rect 250 -2071 256 -1583
rect 273 -2071 279 -1583
rect 250 -2077 279 -2071
rect -279 -2192 -250 -2186
rect -279 -2680 -273 -2192
rect -256 -2680 -250 -2192
rect -279 -2686 -250 -2680
rect 250 -2192 279 -2186
rect 250 -2680 256 -2192
rect 273 -2680 279 -2192
rect 250 -2686 279 -2680
rect -279 -2801 -250 -2795
rect -279 -3289 -273 -2801
rect -256 -3289 -250 -2801
rect -279 -3295 -250 -3289
rect 250 -2801 279 -2795
rect 250 -3289 256 -2801
rect 273 -3289 279 -2801
rect 250 -3295 279 -3289
rect -279 -3410 -250 -3404
rect -279 -3898 -273 -3410
rect -256 -3898 -250 -3410
rect -279 -3904 -250 -3898
rect 250 -3410 279 -3404
rect 250 -3898 256 -3410
rect 273 -3898 279 -3410
rect 250 -3904 279 -3898
rect -279 -4019 -250 -4013
rect -279 -4507 -273 -4019
rect -256 -4507 -250 -4019
rect -279 -4513 -250 -4507
rect 250 -4019 279 -4013
rect 250 -4507 256 -4019
rect 273 -4507 279 -4019
rect 250 -4513 279 -4507
<< ndiffc >>
rect -273 4019 -256 4507
rect 256 4019 273 4507
rect -273 3410 -256 3898
rect 256 3410 273 3898
rect -273 2801 -256 3289
rect 256 2801 273 3289
rect -273 2192 -256 2680
rect 256 2192 273 2680
rect -273 1583 -256 2071
rect 256 1583 273 2071
rect -273 974 -256 1462
rect 256 974 273 1462
rect -273 365 -256 853
rect 256 365 273 853
rect -273 -244 -256 244
rect 256 -244 273 244
rect -273 -853 -256 -365
rect 256 -853 273 -365
rect -273 -1462 -256 -974
rect 256 -1462 273 -974
rect -273 -2071 -256 -1583
rect 256 -2071 273 -1583
rect -273 -2680 -256 -2192
rect 256 -2680 273 -2192
rect -273 -3289 -256 -2801
rect 256 -3289 273 -2801
rect -273 -3898 -256 -3410
rect 256 -3898 273 -3410
rect -273 -4507 -256 -4019
rect 256 -4507 273 -4019
<< poly >>
rect -250 4549 250 4557
rect -250 4532 -242 4549
rect 242 4532 250 4549
rect -250 4513 250 4532
rect -250 3994 250 4013
rect -250 3977 -242 3994
rect 242 3977 250 3994
rect -250 3969 250 3977
rect -250 3940 250 3948
rect -250 3923 -242 3940
rect 242 3923 250 3940
rect -250 3904 250 3923
rect -250 3385 250 3404
rect -250 3368 -242 3385
rect 242 3368 250 3385
rect -250 3360 250 3368
rect -250 3331 250 3339
rect -250 3314 -242 3331
rect 242 3314 250 3331
rect -250 3295 250 3314
rect -250 2776 250 2795
rect -250 2759 -242 2776
rect 242 2759 250 2776
rect -250 2751 250 2759
rect -250 2722 250 2730
rect -250 2705 -242 2722
rect 242 2705 250 2722
rect -250 2686 250 2705
rect -250 2167 250 2186
rect -250 2150 -242 2167
rect 242 2150 250 2167
rect -250 2142 250 2150
rect -250 2113 250 2121
rect -250 2096 -242 2113
rect 242 2096 250 2113
rect -250 2077 250 2096
rect -250 1558 250 1577
rect -250 1541 -242 1558
rect 242 1541 250 1558
rect -250 1533 250 1541
rect -250 1504 250 1512
rect -250 1487 -242 1504
rect 242 1487 250 1504
rect -250 1468 250 1487
rect -250 949 250 968
rect -250 932 -242 949
rect 242 932 250 949
rect -250 924 250 932
rect -250 895 250 903
rect -250 878 -242 895
rect 242 878 250 895
rect -250 859 250 878
rect -250 340 250 359
rect -250 323 -242 340
rect 242 323 250 340
rect -250 315 250 323
rect -250 286 250 294
rect -250 269 -242 286
rect 242 269 250 286
rect -250 250 250 269
rect -250 -269 250 -250
rect -250 -286 -242 -269
rect 242 -286 250 -269
rect -250 -294 250 -286
rect -250 -323 250 -315
rect -250 -340 -242 -323
rect 242 -340 250 -323
rect -250 -359 250 -340
rect -250 -878 250 -859
rect -250 -895 -242 -878
rect 242 -895 250 -878
rect -250 -903 250 -895
rect -250 -932 250 -924
rect -250 -949 -242 -932
rect 242 -949 250 -932
rect -250 -968 250 -949
rect -250 -1487 250 -1468
rect -250 -1504 -242 -1487
rect 242 -1504 250 -1487
rect -250 -1512 250 -1504
rect -250 -1541 250 -1533
rect -250 -1558 -242 -1541
rect 242 -1558 250 -1541
rect -250 -1577 250 -1558
rect -250 -2096 250 -2077
rect -250 -2113 -242 -2096
rect 242 -2113 250 -2096
rect -250 -2121 250 -2113
rect -250 -2150 250 -2142
rect -250 -2167 -242 -2150
rect 242 -2167 250 -2150
rect -250 -2186 250 -2167
rect -250 -2705 250 -2686
rect -250 -2722 -242 -2705
rect 242 -2722 250 -2705
rect -250 -2730 250 -2722
rect -250 -2759 250 -2751
rect -250 -2776 -242 -2759
rect 242 -2776 250 -2759
rect -250 -2795 250 -2776
rect -250 -3314 250 -3295
rect -250 -3331 -242 -3314
rect 242 -3331 250 -3314
rect -250 -3339 250 -3331
rect -250 -3368 250 -3360
rect -250 -3385 -242 -3368
rect 242 -3385 250 -3368
rect -250 -3404 250 -3385
rect -250 -3923 250 -3904
rect -250 -3940 -242 -3923
rect 242 -3940 250 -3923
rect -250 -3948 250 -3940
rect -250 -3977 250 -3969
rect -250 -3994 -242 -3977
rect 242 -3994 250 -3977
rect -250 -4013 250 -3994
rect -250 -4532 250 -4513
rect -250 -4549 -242 -4532
rect 242 -4549 250 -4532
rect -250 -4557 250 -4549
<< polycont >>
rect -242 4532 242 4549
rect -242 3977 242 3994
rect -242 3923 242 3940
rect -242 3368 242 3385
rect -242 3314 242 3331
rect -242 2759 242 2776
rect -242 2705 242 2722
rect -242 2150 242 2167
rect -242 2096 242 2113
rect -242 1541 242 1558
rect -242 1487 242 1504
rect -242 932 242 949
rect -242 878 242 895
rect -242 323 242 340
rect -242 269 242 286
rect -242 -286 242 -269
rect -242 -340 242 -323
rect -242 -895 242 -878
rect -242 -949 242 -932
rect -242 -1504 242 -1487
rect -242 -1558 242 -1541
rect -242 -2113 242 -2096
rect -242 -2167 242 -2150
rect -242 -2722 242 -2705
rect -242 -2776 242 -2759
rect -242 -3331 242 -3314
rect -242 -3385 242 -3368
rect -242 -3940 242 -3923
rect -242 -3994 242 -3977
rect -242 -4549 242 -4532
<< locali >>
rect -250 4532 -242 4549
rect 242 4532 250 4549
rect -273 4507 -256 4515
rect -273 4011 -256 4019
rect 256 4507 273 4515
rect 256 4011 273 4019
rect -250 3977 -242 3994
rect 242 3977 250 3994
rect -250 3923 -242 3940
rect 242 3923 250 3940
rect -273 3898 -256 3906
rect -273 3402 -256 3410
rect 256 3898 273 3906
rect 256 3402 273 3410
rect -250 3368 -242 3385
rect 242 3368 250 3385
rect -250 3314 -242 3331
rect 242 3314 250 3331
rect -273 3289 -256 3297
rect -273 2793 -256 2801
rect 256 3289 273 3297
rect 256 2793 273 2801
rect -250 2759 -242 2776
rect 242 2759 250 2776
rect -250 2705 -242 2722
rect 242 2705 250 2722
rect -273 2680 -256 2688
rect -273 2184 -256 2192
rect 256 2680 273 2688
rect 256 2184 273 2192
rect -250 2150 -242 2167
rect 242 2150 250 2167
rect -250 2096 -242 2113
rect 242 2096 250 2113
rect -273 2071 -256 2079
rect -273 1575 -256 1583
rect 256 2071 273 2079
rect 256 1575 273 1583
rect -250 1541 -242 1558
rect 242 1541 250 1558
rect -250 1487 -242 1504
rect 242 1487 250 1504
rect -273 1462 -256 1470
rect -273 966 -256 974
rect 256 1462 273 1470
rect 256 966 273 974
rect -250 932 -242 949
rect 242 932 250 949
rect -250 878 -242 895
rect 242 878 250 895
rect -273 853 -256 861
rect -273 357 -256 365
rect 256 853 273 861
rect 256 357 273 365
rect -250 323 -242 340
rect 242 323 250 340
rect -250 269 -242 286
rect 242 269 250 286
rect -273 244 -256 252
rect -273 -252 -256 -244
rect 256 244 273 252
rect 256 -252 273 -244
rect -250 -286 -242 -269
rect 242 -286 250 -269
rect -250 -340 -242 -323
rect 242 -340 250 -323
rect -273 -365 -256 -357
rect -273 -861 -256 -853
rect 256 -365 273 -357
rect 256 -861 273 -853
rect -250 -895 -242 -878
rect 242 -895 250 -878
rect -250 -949 -242 -932
rect 242 -949 250 -932
rect -273 -974 -256 -966
rect -273 -1470 -256 -1462
rect 256 -974 273 -966
rect 256 -1470 273 -1462
rect -250 -1504 -242 -1487
rect 242 -1504 250 -1487
rect -250 -1558 -242 -1541
rect 242 -1558 250 -1541
rect -273 -1583 -256 -1575
rect -273 -2079 -256 -2071
rect 256 -1583 273 -1575
rect 256 -2079 273 -2071
rect -250 -2113 -242 -2096
rect 242 -2113 250 -2096
rect -250 -2167 -242 -2150
rect 242 -2167 250 -2150
rect -273 -2192 -256 -2184
rect -273 -2688 -256 -2680
rect 256 -2192 273 -2184
rect 256 -2688 273 -2680
rect -250 -2722 -242 -2705
rect 242 -2722 250 -2705
rect -250 -2776 -242 -2759
rect 242 -2776 250 -2759
rect -273 -2801 -256 -2793
rect -273 -3297 -256 -3289
rect 256 -2801 273 -2793
rect 256 -3297 273 -3289
rect -250 -3331 -242 -3314
rect 242 -3331 250 -3314
rect -250 -3385 -242 -3368
rect 242 -3385 250 -3368
rect -273 -3410 -256 -3402
rect -273 -3906 -256 -3898
rect 256 -3410 273 -3402
rect 256 -3906 273 -3898
rect -250 -3940 -242 -3923
rect 242 -3940 250 -3923
rect -250 -3994 -242 -3977
rect 242 -3994 250 -3977
rect -273 -4019 -256 -4011
rect -273 -4515 -256 -4507
rect 256 -4019 273 -4011
rect 256 -4515 273 -4507
rect -250 -4549 -242 -4532
rect 242 -4549 250 -4532
<< viali >>
rect -242 4532 242 4549
rect -273 4019 -256 4507
rect 256 4019 273 4507
rect -242 3977 242 3994
rect -242 3923 242 3940
rect -273 3410 -256 3898
rect 256 3410 273 3898
rect -242 3368 242 3385
rect -242 3314 242 3331
rect -273 2801 -256 3289
rect 256 2801 273 3289
rect -242 2759 242 2776
rect -242 2705 242 2722
rect -273 2192 -256 2680
rect 256 2192 273 2680
rect -242 2150 242 2167
rect -242 2096 242 2113
rect -273 1583 -256 2071
rect 256 1583 273 2071
rect -242 1541 242 1558
rect -242 1487 242 1504
rect -273 974 -256 1462
rect 256 974 273 1462
rect -242 932 242 949
rect -242 878 242 895
rect -273 365 -256 853
rect 256 365 273 853
rect -242 323 242 340
rect -242 269 242 286
rect -273 -244 -256 244
rect 256 -244 273 244
rect -242 -286 242 -269
rect -242 -340 242 -323
rect -273 -853 -256 -365
rect 256 -853 273 -365
rect -242 -895 242 -878
rect -242 -949 242 -932
rect -273 -1462 -256 -974
rect 256 -1462 273 -974
rect -242 -1504 242 -1487
rect -242 -1558 242 -1541
rect -273 -2071 -256 -1583
rect 256 -2071 273 -1583
rect -242 -2113 242 -2096
rect -242 -2167 242 -2150
rect -273 -2680 -256 -2192
rect 256 -2680 273 -2192
rect -242 -2722 242 -2705
rect -242 -2776 242 -2759
rect -273 -3289 -256 -2801
rect 256 -3289 273 -2801
rect -242 -3331 242 -3314
rect -242 -3385 242 -3368
rect -273 -3898 -256 -3410
rect 256 -3898 273 -3410
rect -242 -3940 242 -3923
rect -242 -3994 242 -3977
rect -273 -4507 -256 -4019
rect 256 -4507 273 -4019
rect -242 -4549 242 -4532
<< metal1 >>
rect -248 4549 248 4552
rect -248 4532 -242 4549
rect 242 4532 248 4549
rect -248 4529 248 4532
rect -276 4507 -253 4513
rect -276 4019 -273 4507
rect -256 4019 -253 4507
rect -276 4013 -253 4019
rect 253 4507 276 4513
rect 253 4019 256 4507
rect 273 4019 276 4507
rect 253 4013 276 4019
rect -248 3994 248 3997
rect -248 3977 -242 3994
rect 242 3977 248 3994
rect -248 3974 248 3977
rect -248 3940 248 3943
rect -248 3923 -242 3940
rect 242 3923 248 3940
rect -248 3920 248 3923
rect -276 3898 -253 3904
rect -276 3410 -273 3898
rect -256 3410 -253 3898
rect -276 3404 -253 3410
rect 253 3898 276 3904
rect 253 3410 256 3898
rect 273 3410 276 3898
rect 253 3404 276 3410
rect -248 3385 248 3388
rect -248 3368 -242 3385
rect 242 3368 248 3385
rect -248 3365 248 3368
rect -248 3331 248 3334
rect -248 3314 -242 3331
rect 242 3314 248 3331
rect -248 3311 248 3314
rect -276 3289 -253 3295
rect -276 2801 -273 3289
rect -256 2801 -253 3289
rect -276 2795 -253 2801
rect 253 3289 276 3295
rect 253 2801 256 3289
rect 273 2801 276 3289
rect 253 2795 276 2801
rect -248 2776 248 2779
rect -248 2759 -242 2776
rect 242 2759 248 2776
rect -248 2756 248 2759
rect -248 2722 248 2725
rect -248 2705 -242 2722
rect 242 2705 248 2722
rect -248 2702 248 2705
rect -276 2680 -253 2686
rect -276 2192 -273 2680
rect -256 2192 -253 2680
rect -276 2186 -253 2192
rect 253 2680 276 2686
rect 253 2192 256 2680
rect 273 2192 276 2680
rect 253 2186 276 2192
rect -248 2167 248 2170
rect -248 2150 -242 2167
rect 242 2150 248 2167
rect -248 2147 248 2150
rect -248 2113 248 2116
rect -248 2096 -242 2113
rect 242 2096 248 2113
rect -248 2093 248 2096
rect -276 2071 -253 2077
rect -276 1583 -273 2071
rect -256 1583 -253 2071
rect -276 1577 -253 1583
rect 253 2071 276 2077
rect 253 1583 256 2071
rect 273 1583 276 2071
rect 253 1577 276 1583
rect -248 1558 248 1561
rect -248 1541 -242 1558
rect 242 1541 248 1558
rect -248 1538 248 1541
rect -248 1504 248 1507
rect -248 1487 -242 1504
rect 242 1487 248 1504
rect -248 1484 248 1487
rect -276 1462 -253 1468
rect -276 974 -273 1462
rect -256 974 -253 1462
rect -276 968 -253 974
rect 253 1462 276 1468
rect 253 974 256 1462
rect 273 974 276 1462
rect 253 968 276 974
rect -248 949 248 952
rect -248 932 -242 949
rect 242 932 248 949
rect -248 929 248 932
rect -248 895 248 898
rect -248 878 -242 895
rect 242 878 248 895
rect -248 875 248 878
rect -276 853 -253 859
rect -276 365 -273 853
rect -256 365 -253 853
rect -276 359 -253 365
rect 253 853 276 859
rect 253 365 256 853
rect 273 365 276 853
rect 253 359 276 365
rect -248 340 248 343
rect -248 323 -242 340
rect 242 323 248 340
rect -248 320 248 323
rect -248 286 248 289
rect -248 269 -242 286
rect 242 269 248 286
rect -248 266 248 269
rect -276 244 -253 250
rect -276 -244 -273 244
rect -256 -244 -253 244
rect -276 -250 -253 -244
rect 253 244 276 250
rect 253 -244 256 244
rect 273 -244 276 244
rect 253 -250 276 -244
rect -248 -269 248 -266
rect -248 -286 -242 -269
rect 242 -286 248 -269
rect -248 -289 248 -286
rect -248 -323 248 -320
rect -248 -340 -242 -323
rect 242 -340 248 -323
rect -248 -343 248 -340
rect -276 -365 -253 -359
rect -276 -853 -273 -365
rect -256 -853 -253 -365
rect -276 -859 -253 -853
rect 253 -365 276 -359
rect 253 -853 256 -365
rect 273 -853 276 -365
rect 253 -859 276 -853
rect -248 -878 248 -875
rect -248 -895 -242 -878
rect 242 -895 248 -878
rect -248 -898 248 -895
rect -248 -932 248 -929
rect -248 -949 -242 -932
rect 242 -949 248 -932
rect -248 -952 248 -949
rect -276 -974 -253 -968
rect -276 -1462 -273 -974
rect -256 -1462 -253 -974
rect -276 -1468 -253 -1462
rect 253 -974 276 -968
rect 253 -1462 256 -974
rect 273 -1462 276 -974
rect 253 -1468 276 -1462
rect -248 -1487 248 -1484
rect -248 -1504 -242 -1487
rect 242 -1504 248 -1487
rect -248 -1507 248 -1504
rect -248 -1541 248 -1538
rect -248 -1558 -242 -1541
rect 242 -1558 248 -1541
rect -248 -1561 248 -1558
rect -276 -1583 -253 -1577
rect -276 -2071 -273 -1583
rect -256 -2071 -253 -1583
rect -276 -2077 -253 -2071
rect 253 -1583 276 -1577
rect 253 -2071 256 -1583
rect 273 -2071 276 -1583
rect 253 -2077 276 -2071
rect -248 -2096 248 -2093
rect -248 -2113 -242 -2096
rect 242 -2113 248 -2096
rect -248 -2116 248 -2113
rect -248 -2150 248 -2147
rect -248 -2167 -242 -2150
rect 242 -2167 248 -2150
rect -248 -2170 248 -2167
rect -276 -2192 -253 -2186
rect -276 -2680 -273 -2192
rect -256 -2680 -253 -2192
rect -276 -2686 -253 -2680
rect 253 -2192 276 -2186
rect 253 -2680 256 -2192
rect 273 -2680 276 -2192
rect 253 -2686 276 -2680
rect -248 -2705 248 -2702
rect -248 -2722 -242 -2705
rect 242 -2722 248 -2705
rect -248 -2725 248 -2722
rect -248 -2759 248 -2756
rect -248 -2776 -242 -2759
rect 242 -2776 248 -2759
rect -248 -2779 248 -2776
rect -276 -2801 -253 -2795
rect -276 -3289 -273 -2801
rect -256 -3289 -253 -2801
rect -276 -3295 -253 -3289
rect 253 -2801 276 -2795
rect 253 -3289 256 -2801
rect 273 -3289 276 -2801
rect 253 -3295 276 -3289
rect -248 -3314 248 -3311
rect -248 -3331 -242 -3314
rect 242 -3331 248 -3314
rect -248 -3334 248 -3331
rect -248 -3368 248 -3365
rect -248 -3385 -242 -3368
rect 242 -3385 248 -3368
rect -248 -3388 248 -3385
rect -276 -3410 -253 -3404
rect -276 -3898 -273 -3410
rect -256 -3898 -253 -3410
rect -276 -3904 -253 -3898
rect 253 -3410 276 -3404
rect 253 -3898 256 -3410
rect 273 -3898 276 -3410
rect 253 -3904 276 -3898
rect -248 -3923 248 -3920
rect -248 -3940 -242 -3923
rect 242 -3940 248 -3923
rect -248 -3943 248 -3940
rect -248 -3977 248 -3974
rect -248 -3994 -242 -3977
rect 242 -3994 248 -3977
rect -248 -3997 248 -3994
rect -276 -4019 -253 -4013
rect -276 -4507 -273 -4019
rect -256 -4507 -253 -4019
rect -276 -4513 -253 -4507
rect 253 -4019 276 -4013
rect 253 -4507 256 -4019
rect 273 -4507 276 -4019
rect 253 -4513 276 -4507
rect -248 -4532 248 -4529
rect -248 -4549 -242 -4532
rect 242 -4549 248 -4532
rect -248 -4552 248 -4549
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 5.0 l 5.0 m 15 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
