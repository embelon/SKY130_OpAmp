magic
tech sky130A
magscale 1 2
timestamp 1695663670
<< error_p >>
rect -1594 61818 1594 62036
rect -1594 60582 1594 60800
rect -1594 59346 1594 59564
rect -1594 58110 1594 58328
rect -1594 56874 1594 57092
rect -1594 55638 1594 55856
rect -1594 54402 1594 54620
rect -1594 53166 1594 53384
rect -1594 51930 1594 52148
rect -1594 50694 1594 50912
rect -1594 49458 1594 49676
rect -1594 48222 1594 48440
rect -1594 46986 1594 47204
rect -1594 45750 1594 45968
rect -1594 44514 1594 44732
rect -1594 43278 1594 43496
rect -1594 42042 1594 42260
rect -1594 40806 1594 41024
rect -1594 39570 1594 39788
rect -1594 38334 1594 38552
rect -1594 37098 1594 37316
rect -1594 35862 1594 36080
rect -1594 34626 1594 34844
rect -1594 33390 1594 33608
rect -1594 32154 1594 32372
rect -1594 30918 1594 31136
rect -1594 29682 1594 29900
rect -1594 28446 1594 28664
rect -1594 27210 1594 27428
rect -1594 25974 1594 26192
rect -1594 24738 1594 24956
rect -1594 23502 1594 23720
rect -1594 22266 1594 22484
rect -1594 21030 1594 21248
rect -1594 19794 1594 20012
rect -1594 18558 1594 18776
rect -1594 17322 1594 17540
rect -1594 16086 1594 16304
rect -1594 14850 1594 15068
rect -1594 13614 1594 13832
rect -1594 12378 1594 12596
rect -1594 11142 1594 11360
rect -1594 9906 1594 10124
rect -1594 8670 1594 8888
rect -1594 7434 1594 7652
rect -1594 6198 1594 6416
rect -1594 4962 1594 5180
rect -1594 3726 1594 3944
rect -1594 2490 1594 2708
rect -1594 1254 1594 1472
rect -1594 18 1594 236
rect -1594 -1218 1594 -1000
rect -1594 -2454 1594 -2236
rect -1594 -3690 1594 -3472
rect -1594 -4926 1594 -4708
rect -1594 -6162 1594 -5944
rect -1594 -7398 1594 -7180
rect -1594 -8634 1594 -8416
rect -1594 -9870 1594 -9652
rect -1594 -11106 1594 -10888
rect -1594 -12342 1594 -12124
rect -1594 -13578 1594 -13360
rect -1594 -14814 1594 -14596
rect -1594 -16050 1594 -15832
rect -1594 -17286 1594 -17068
rect -1594 -18522 1594 -18304
rect -1594 -19758 1594 -19540
rect -1594 -20994 1594 -20776
rect -1594 -22230 1594 -22012
rect -1594 -23466 1594 -23248
rect -1594 -24702 1594 -24484
rect -1594 -25938 1594 -25720
rect -1594 -27174 1594 -26956
rect -1594 -28410 1594 -28192
rect -1594 -29646 1594 -29428
rect -1594 -30882 1594 -30664
rect -1594 -32118 1594 -31900
rect -1594 -33354 1594 -33136
rect -1594 -34590 1594 -34372
rect -1594 -35826 1594 -35608
rect -1594 -37062 1594 -36844
rect -1594 -38298 1594 -38080
rect -1594 -39534 1594 -39316
rect -1594 -40770 1594 -40552
rect -1594 -42006 1594 -41788
rect -1594 -43242 1594 -43024
rect -1594 -44478 1594 -44260
rect -1594 -45714 1594 -45496
rect -1594 -46950 1594 -46732
rect -1594 -48186 1594 -47968
rect -1594 -49422 1594 -49204
rect -1594 -50658 1594 -50440
rect -1594 -51894 1594 -51676
rect -1594 -53130 1594 -52912
rect -1594 -54366 1594 -54148
rect -1594 -55602 1594 -55384
rect -1594 -56838 1594 -56620
rect -1594 -58074 1594 -57856
rect -1594 -59310 1594 -59092
rect -1594 -60546 1594 -60328
rect -1594 -61782 1594 -61564
<< nwell >>
rect -1594 61818 1594 63018
rect -1594 60582 1594 61782
rect -1594 59346 1594 60546
rect -1594 58110 1594 59310
rect -1594 56874 1594 58074
rect -1594 55638 1594 56838
rect -1594 54402 1594 55602
rect -1594 53166 1594 54366
rect -1594 51930 1594 53130
rect -1594 50694 1594 51894
rect -1594 49458 1594 50658
rect -1594 48222 1594 49422
rect -1594 46986 1594 48186
rect -1594 45750 1594 46950
rect -1594 44514 1594 45714
rect -1594 43278 1594 44478
rect -1594 42042 1594 43242
rect -1594 40806 1594 42006
rect -1594 39570 1594 40770
rect -1594 38334 1594 39534
rect -1594 37098 1594 38298
rect -1594 35862 1594 37062
rect -1594 34626 1594 35826
rect -1594 33390 1594 34590
rect -1594 32154 1594 33354
rect -1594 30918 1594 32118
rect -1594 29682 1594 30882
rect -1594 28446 1594 29646
rect -1594 27210 1594 28410
rect -1594 25974 1594 27174
rect -1594 24738 1594 25938
rect -1594 23502 1594 24702
rect -1594 22266 1594 23466
rect -1594 21030 1594 22230
rect -1594 19794 1594 20994
rect -1594 18558 1594 19758
rect -1594 17322 1594 18522
rect -1594 16086 1594 17286
rect -1594 14850 1594 16050
rect -1594 13614 1594 14814
rect -1594 12378 1594 13578
rect -1594 11142 1594 12342
rect -1594 9906 1594 11106
rect -1594 8670 1594 9870
rect -1594 7434 1594 8634
rect -1594 6198 1594 7398
rect -1594 4962 1594 6162
rect -1594 3726 1594 4926
rect -1594 2490 1594 3690
rect -1594 1254 1594 2454
rect -1594 18 1594 1218
rect -1594 -1218 1594 -18
rect -1594 -2454 1594 -1254
rect -1594 -3690 1594 -2490
rect -1594 -4926 1594 -3726
rect -1594 -6162 1594 -4962
rect -1594 -7398 1594 -6198
rect -1594 -8634 1594 -7434
rect -1594 -9870 1594 -8670
rect -1594 -11106 1594 -9906
rect -1594 -12342 1594 -11142
rect -1594 -13578 1594 -12378
rect -1594 -14814 1594 -13614
rect -1594 -16050 1594 -14850
rect -1594 -17286 1594 -16086
rect -1594 -18522 1594 -17322
rect -1594 -19758 1594 -18558
rect -1594 -20994 1594 -19794
rect -1594 -22230 1594 -21030
rect -1594 -23466 1594 -22266
rect -1594 -24702 1594 -23502
rect -1594 -25938 1594 -24738
rect -1594 -27174 1594 -25974
rect -1594 -28410 1594 -27210
rect -1594 -29646 1594 -28446
rect -1594 -30882 1594 -29682
rect -1594 -32118 1594 -30918
rect -1594 -33354 1594 -32154
rect -1594 -34590 1594 -33390
rect -1594 -35826 1594 -34626
rect -1594 -37062 1594 -35862
rect -1594 -38298 1594 -37098
rect -1594 -39534 1594 -38334
rect -1594 -40770 1594 -39570
rect -1594 -42006 1594 -40806
rect -1594 -43242 1594 -42042
rect -1594 -44478 1594 -43278
rect -1594 -45714 1594 -44514
rect -1594 -46950 1594 -45750
rect -1594 -48186 1594 -46986
rect -1594 -49422 1594 -48222
rect -1594 -50658 1594 -49458
rect -1594 -51894 1594 -50694
rect -1594 -53130 1594 -51930
rect -1594 -54366 1594 -53166
rect -1594 -55602 1594 -54402
rect -1594 -56838 1594 -55638
rect -1594 -58074 1594 -56874
rect -1594 -59310 1594 -58110
rect -1594 -60546 1594 -59346
rect -1594 -61782 1594 -60582
rect -1594 -63018 1594 -61818
<< pmos >>
rect -1500 61918 1500 62918
rect -1500 60682 1500 61682
rect -1500 59446 1500 60446
rect -1500 58210 1500 59210
rect -1500 56974 1500 57974
rect -1500 55738 1500 56738
rect -1500 54502 1500 55502
rect -1500 53266 1500 54266
rect -1500 52030 1500 53030
rect -1500 50794 1500 51794
rect -1500 49558 1500 50558
rect -1500 48322 1500 49322
rect -1500 47086 1500 48086
rect -1500 45850 1500 46850
rect -1500 44614 1500 45614
rect -1500 43378 1500 44378
rect -1500 42142 1500 43142
rect -1500 40906 1500 41906
rect -1500 39670 1500 40670
rect -1500 38434 1500 39434
rect -1500 37198 1500 38198
rect -1500 35962 1500 36962
rect -1500 34726 1500 35726
rect -1500 33490 1500 34490
rect -1500 32254 1500 33254
rect -1500 31018 1500 32018
rect -1500 29782 1500 30782
rect -1500 28546 1500 29546
rect -1500 27310 1500 28310
rect -1500 26074 1500 27074
rect -1500 24838 1500 25838
rect -1500 23602 1500 24602
rect -1500 22366 1500 23366
rect -1500 21130 1500 22130
rect -1500 19894 1500 20894
rect -1500 18658 1500 19658
rect -1500 17422 1500 18422
rect -1500 16186 1500 17186
rect -1500 14950 1500 15950
rect -1500 13714 1500 14714
rect -1500 12478 1500 13478
rect -1500 11242 1500 12242
rect -1500 10006 1500 11006
rect -1500 8770 1500 9770
rect -1500 7534 1500 8534
rect -1500 6298 1500 7298
rect -1500 5062 1500 6062
rect -1500 3826 1500 4826
rect -1500 2590 1500 3590
rect -1500 1354 1500 2354
rect -1500 118 1500 1118
rect -1500 -1118 1500 -118
rect -1500 -2354 1500 -1354
rect -1500 -3590 1500 -2590
rect -1500 -4826 1500 -3826
rect -1500 -6062 1500 -5062
rect -1500 -7298 1500 -6298
rect -1500 -8534 1500 -7534
rect -1500 -9770 1500 -8770
rect -1500 -11006 1500 -10006
rect -1500 -12242 1500 -11242
rect -1500 -13478 1500 -12478
rect -1500 -14714 1500 -13714
rect -1500 -15950 1500 -14950
rect -1500 -17186 1500 -16186
rect -1500 -18422 1500 -17422
rect -1500 -19658 1500 -18658
rect -1500 -20894 1500 -19894
rect -1500 -22130 1500 -21130
rect -1500 -23366 1500 -22366
rect -1500 -24602 1500 -23602
rect -1500 -25838 1500 -24838
rect -1500 -27074 1500 -26074
rect -1500 -28310 1500 -27310
rect -1500 -29546 1500 -28546
rect -1500 -30782 1500 -29782
rect -1500 -32018 1500 -31018
rect -1500 -33254 1500 -32254
rect -1500 -34490 1500 -33490
rect -1500 -35726 1500 -34726
rect -1500 -36962 1500 -35962
rect -1500 -38198 1500 -37198
rect -1500 -39434 1500 -38434
rect -1500 -40670 1500 -39670
rect -1500 -41906 1500 -40906
rect -1500 -43142 1500 -42142
rect -1500 -44378 1500 -43378
rect -1500 -45614 1500 -44614
rect -1500 -46850 1500 -45850
rect -1500 -48086 1500 -47086
rect -1500 -49322 1500 -48322
rect -1500 -50558 1500 -49558
rect -1500 -51794 1500 -50794
rect -1500 -53030 1500 -52030
rect -1500 -54266 1500 -53266
rect -1500 -55502 1500 -54502
rect -1500 -56738 1500 -55738
rect -1500 -57974 1500 -56974
rect -1500 -59210 1500 -58210
rect -1500 -60446 1500 -59446
rect -1500 -61682 1500 -60682
rect -1500 -62918 1500 -61918
<< pdiff >>
rect -1558 62906 -1500 62918
rect -1558 61930 -1546 62906
rect -1512 61930 -1500 62906
rect -1558 61918 -1500 61930
rect 1500 62906 1558 62918
rect 1500 61930 1512 62906
rect 1546 61930 1558 62906
rect 1500 61918 1558 61930
rect -1558 61670 -1500 61682
rect -1558 60694 -1546 61670
rect -1512 60694 -1500 61670
rect -1558 60682 -1500 60694
rect 1500 61670 1558 61682
rect 1500 60694 1512 61670
rect 1546 60694 1558 61670
rect 1500 60682 1558 60694
rect -1558 60434 -1500 60446
rect -1558 59458 -1546 60434
rect -1512 59458 -1500 60434
rect -1558 59446 -1500 59458
rect 1500 60434 1558 60446
rect 1500 59458 1512 60434
rect 1546 59458 1558 60434
rect 1500 59446 1558 59458
rect -1558 59198 -1500 59210
rect -1558 58222 -1546 59198
rect -1512 58222 -1500 59198
rect -1558 58210 -1500 58222
rect 1500 59198 1558 59210
rect 1500 58222 1512 59198
rect 1546 58222 1558 59198
rect 1500 58210 1558 58222
rect -1558 57962 -1500 57974
rect -1558 56986 -1546 57962
rect -1512 56986 -1500 57962
rect -1558 56974 -1500 56986
rect 1500 57962 1558 57974
rect 1500 56986 1512 57962
rect 1546 56986 1558 57962
rect 1500 56974 1558 56986
rect -1558 56726 -1500 56738
rect -1558 55750 -1546 56726
rect -1512 55750 -1500 56726
rect -1558 55738 -1500 55750
rect 1500 56726 1558 56738
rect 1500 55750 1512 56726
rect 1546 55750 1558 56726
rect 1500 55738 1558 55750
rect -1558 55490 -1500 55502
rect -1558 54514 -1546 55490
rect -1512 54514 -1500 55490
rect -1558 54502 -1500 54514
rect 1500 55490 1558 55502
rect 1500 54514 1512 55490
rect 1546 54514 1558 55490
rect 1500 54502 1558 54514
rect -1558 54254 -1500 54266
rect -1558 53278 -1546 54254
rect -1512 53278 -1500 54254
rect -1558 53266 -1500 53278
rect 1500 54254 1558 54266
rect 1500 53278 1512 54254
rect 1546 53278 1558 54254
rect 1500 53266 1558 53278
rect -1558 53018 -1500 53030
rect -1558 52042 -1546 53018
rect -1512 52042 -1500 53018
rect -1558 52030 -1500 52042
rect 1500 53018 1558 53030
rect 1500 52042 1512 53018
rect 1546 52042 1558 53018
rect 1500 52030 1558 52042
rect -1558 51782 -1500 51794
rect -1558 50806 -1546 51782
rect -1512 50806 -1500 51782
rect -1558 50794 -1500 50806
rect 1500 51782 1558 51794
rect 1500 50806 1512 51782
rect 1546 50806 1558 51782
rect 1500 50794 1558 50806
rect -1558 50546 -1500 50558
rect -1558 49570 -1546 50546
rect -1512 49570 -1500 50546
rect -1558 49558 -1500 49570
rect 1500 50546 1558 50558
rect 1500 49570 1512 50546
rect 1546 49570 1558 50546
rect 1500 49558 1558 49570
rect -1558 49310 -1500 49322
rect -1558 48334 -1546 49310
rect -1512 48334 -1500 49310
rect -1558 48322 -1500 48334
rect 1500 49310 1558 49322
rect 1500 48334 1512 49310
rect 1546 48334 1558 49310
rect 1500 48322 1558 48334
rect -1558 48074 -1500 48086
rect -1558 47098 -1546 48074
rect -1512 47098 -1500 48074
rect -1558 47086 -1500 47098
rect 1500 48074 1558 48086
rect 1500 47098 1512 48074
rect 1546 47098 1558 48074
rect 1500 47086 1558 47098
rect -1558 46838 -1500 46850
rect -1558 45862 -1546 46838
rect -1512 45862 -1500 46838
rect -1558 45850 -1500 45862
rect 1500 46838 1558 46850
rect 1500 45862 1512 46838
rect 1546 45862 1558 46838
rect 1500 45850 1558 45862
rect -1558 45602 -1500 45614
rect -1558 44626 -1546 45602
rect -1512 44626 -1500 45602
rect -1558 44614 -1500 44626
rect 1500 45602 1558 45614
rect 1500 44626 1512 45602
rect 1546 44626 1558 45602
rect 1500 44614 1558 44626
rect -1558 44366 -1500 44378
rect -1558 43390 -1546 44366
rect -1512 43390 -1500 44366
rect -1558 43378 -1500 43390
rect 1500 44366 1558 44378
rect 1500 43390 1512 44366
rect 1546 43390 1558 44366
rect 1500 43378 1558 43390
rect -1558 43130 -1500 43142
rect -1558 42154 -1546 43130
rect -1512 42154 -1500 43130
rect -1558 42142 -1500 42154
rect 1500 43130 1558 43142
rect 1500 42154 1512 43130
rect 1546 42154 1558 43130
rect 1500 42142 1558 42154
rect -1558 41894 -1500 41906
rect -1558 40918 -1546 41894
rect -1512 40918 -1500 41894
rect -1558 40906 -1500 40918
rect 1500 41894 1558 41906
rect 1500 40918 1512 41894
rect 1546 40918 1558 41894
rect 1500 40906 1558 40918
rect -1558 40658 -1500 40670
rect -1558 39682 -1546 40658
rect -1512 39682 -1500 40658
rect -1558 39670 -1500 39682
rect 1500 40658 1558 40670
rect 1500 39682 1512 40658
rect 1546 39682 1558 40658
rect 1500 39670 1558 39682
rect -1558 39422 -1500 39434
rect -1558 38446 -1546 39422
rect -1512 38446 -1500 39422
rect -1558 38434 -1500 38446
rect 1500 39422 1558 39434
rect 1500 38446 1512 39422
rect 1546 38446 1558 39422
rect 1500 38434 1558 38446
rect -1558 38186 -1500 38198
rect -1558 37210 -1546 38186
rect -1512 37210 -1500 38186
rect -1558 37198 -1500 37210
rect 1500 38186 1558 38198
rect 1500 37210 1512 38186
rect 1546 37210 1558 38186
rect 1500 37198 1558 37210
rect -1558 36950 -1500 36962
rect -1558 35974 -1546 36950
rect -1512 35974 -1500 36950
rect -1558 35962 -1500 35974
rect 1500 36950 1558 36962
rect 1500 35974 1512 36950
rect 1546 35974 1558 36950
rect 1500 35962 1558 35974
rect -1558 35714 -1500 35726
rect -1558 34738 -1546 35714
rect -1512 34738 -1500 35714
rect -1558 34726 -1500 34738
rect 1500 35714 1558 35726
rect 1500 34738 1512 35714
rect 1546 34738 1558 35714
rect 1500 34726 1558 34738
rect -1558 34478 -1500 34490
rect -1558 33502 -1546 34478
rect -1512 33502 -1500 34478
rect -1558 33490 -1500 33502
rect 1500 34478 1558 34490
rect 1500 33502 1512 34478
rect 1546 33502 1558 34478
rect 1500 33490 1558 33502
rect -1558 33242 -1500 33254
rect -1558 32266 -1546 33242
rect -1512 32266 -1500 33242
rect -1558 32254 -1500 32266
rect 1500 33242 1558 33254
rect 1500 32266 1512 33242
rect 1546 32266 1558 33242
rect 1500 32254 1558 32266
rect -1558 32006 -1500 32018
rect -1558 31030 -1546 32006
rect -1512 31030 -1500 32006
rect -1558 31018 -1500 31030
rect 1500 32006 1558 32018
rect 1500 31030 1512 32006
rect 1546 31030 1558 32006
rect 1500 31018 1558 31030
rect -1558 30770 -1500 30782
rect -1558 29794 -1546 30770
rect -1512 29794 -1500 30770
rect -1558 29782 -1500 29794
rect 1500 30770 1558 30782
rect 1500 29794 1512 30770
rect 1546 29794 1558 30770
rect 1500 29782 1558 29794
rect -1558 29534 -1500 29546
rect -1558 28558 -1546 29534
rect -1512 28558 -1500 29534
rect -1558 28546 -1500 28558
rect 1500 29534 1558 29546
rect 1500 28558 1512 29534
rect 1546 28558 1558 29534
rect 1500 28546 1558 28558
rect -1558 28298 -1500 28310
rect -1558 27322 -1546 28298
rect -1512 27322 -1500 28298
rect -1558 27310 -1500 27322
rect 1500 28298 1558 28310
rect 1500 27322 1512 28298
rect 1546 27322 1558 28298
rect 1500 27310 1558 27322
rect -1558 27062 -1500 27074
rect -1558 26086 -1546 27062
rect -1512 26086 -1500 27062
rect -1558 26074 -1500 26086
rect 1500 27062 1558 27074
rect 1500 26086 1512 27062
rect 1546 26086 1558 27062
rect 1500 26074 1558 26086
rect -1558 25826 -1500 25838
rect -1558 24850 -1546 25826
rect -1512 24850 -1500 25826
rect -1558 24838 -1500 24850
rect 1500 25826 1558 25838
rect 1500 24850 1512 25826
rect 1546 24850 1558 25826
rect 1500 24838 1558 24850
rect -1558 24590 -1500 24602
rect -1558 23614 -1546 24590
rect -1512 23614 -1500 24590
rect -1558 23602 -1500 23614
rect 1500 24590 1558 24602
rect 1500 23614 1512 24590
rect 1546 23614 1558 24590
rect 1500 23602 1558 23614
rect -1558 23354 -1500 23366
rect -1558 22378 -1546 23354
rect -1512 22378 -1500 23354
rect -1558 22366 -1500 22378
rect 1500 23354 1558 23366
rect 1500 22378 1512 23354
rect 1546 22378 1558 23354
rect 1500 22366 1558 22378
rect -1558 22118 -1500 22130
rect -1558 21142 -1546 22118
rect -1512 21142 -1500 22118
rect -1558 21130 -1500 21142
rect 1500 22118 1558 22130
rect 1500 21142 1512 22118
rect 1546 21142 1558 22118
rect 1500 21130 1558 21142
rect -1558 20882 -1500 20894
rect -1558 19906 -1546 20882
rect -1512 19906 -1500 20882
rect -1558 19894 -1500 19906
rect 1500 20882 1558 20894
rect 1500 19906 1512 20882
rect 1546 19906 1558 20882
rect 1500 19894 1558 19906
rect -1558 19646 -1500 19658
rect -1558 18670 -1546 19646
rect -1512 18670 -1500 19646
rect -1558 18658 -1500 18670
rect 1500 19646 1558 19658
rect 1500 18670 1512 19646
rect 1546 18670 1558 19646
rect 1500 18658 1558 18670
rect -1558 18410 -1500 18422
rect -1558 17434 -1546 18410
rect -1512 17434 -1500 18410
rect -1558 17422 -1500 17434
rect 1500 18410 1558 18422
rect 1500 17434 1512 18410
rect 1546 17434 1558 18410
rect 1500 17422 1558 17434
rect -1558 17174 -1500 17186
rect -1558 16198 -1546 17174
rect -1512 16198 -1500 17174
rect -1558 16186 -1500 16198
rect 1500 17174 1558 17186
rect 1500 16198 1512 17174
rect 1546 16198 1558 17174
rect 1500 16186 1558 16198
rect -1558 15938 -1500 15950
rect -1558 14962 -1546 15938
rect -1512 14962 -1500 15938
rect -1558 14950 -1500 14962
rect 1500 15938 1558 15950
rect 1500 14962 1512 15938
rect 1546 14962 1558 15938
rect 1500 14950 1558 14962
rect -1558 14702 -1500 14714
rect -1558 13726 -1546 14702
rect -1512 13726 -1500 14702
rect -1558 13714 -1500 13726
rect 1500 14702 1558 14714
rect 1500 13726 1512 14702
rect 1546 13726 1558 14702
rect 1500 13714 1558 13726
rect -1558 13466 -1500 13478
rect -1558 12490 -1546 13466
rect -1512 12490 -1500 13466
rect -1558 12478 -1500 12490
rect 1500 13466 1558 13478
rect 1500 12490 1512 13466
rect 1546 12490 1558 13466
rect 1500 12478 1558 12490
rect -1558 12230 -1500 12242
rect -1558 11254 -1546 12230
rect -1512 11254 -1500 12230
rect -1558 11242 -1500 11254
rect 1500 12230 1558 12242
rect 1500 11254 1512 12230
rect 1546 11254 1558 12230
rect 1500 11242 1558 11254
rect -1558 10994 -1500 11006
rect -1558 10018 -1546 10994
rect -1512 10018 -1500 10994
rect -1558 10006 -1500 10018
rect 1500 10994 1558 11006
rect 1500 10018 1512 10994
rect 1546 10018 1558 10994
rect 1500 10006 1558 10018
rect -1558 9758 -1500 9770
rect -1558 8782 -1546 9758
rect -1512 8782 -1500 9758
rect -1558 8770 -1500 8782
rect 1500 9758 1558 9770
rect 1500 8782 1512 9758
rect 1546 8782 1558 9758
rect 1500 8770 1558 8782
rect -1558 8522 -1500 8534
rect -1558 7546 -1546 8522
rect -1512 7546 -1500 8522
rect -1558 7534 -1500 7546
rect 1500 8522 1558 8534
rect 1500 7546 1512 8522
rect 1546 7546 1558 8522
rect 1500 7534 1558 7546
rect -1558 7286 -1500 7298
rect -1558 6310 -1546 7286
rect -1512 6310 -1500 7286
rect -1558 6298 -1500 6310
rect 1500 7286 1558 7298
rect 1500 6310 1512 7286
rect 1546 6310 1558 7286
rect 1500 6298 1558 6310
rect -1558 6050 -1500 6062
rect -1558 5074 -1546 6050
rect -1512 5074 -1500 6050
rect -1558 5062 -1500 5074
rect 1500 6050 1558 6062
rect 1500 5074 1512 6050
rect 1546 5074 1558 6050
rect 1500 5062 1558 5074
rect -1558 4814 -1500 4826
rect -1558 3838 -1546 4814
rect -1512 3838 -1500 4814
rect -1558 3826 -1500 3838
rect 1500 4814 1558 4826
rect 1500 3838 1512 4814
rect 1546 3838 1558 4814
rect 1500 3826 1558 3838
rect -1558 3578 -1500 3590
rect -1558 2602 -1546 3578
rect -1512 2602 -1500 3578
rect -1558 2590 -1500 2602
rect 1500 3578 1558 3590
rect 1500 2602 1512 3578
rect 1546 2602 1558 3578
rect 1500 2590 1558 2602
rect -1558 2342 -1500 2354
rect -1558 1366 -1546 2342
rect -1512 1366 -1500 2342
rect -1558 1354 -1500 1366
rect 1500 2342 1558 2354
rect 1500 1366 1512 2342
rect 1546 1366 1558 2342
rect 1500 1354 1558 1366
rect -1558 1106 -1500 1118
rect -1558 130 -1546 1106
rect -1512 130 -1500 1106
rect -1558 118 -1500 130
rect 1500 1106 1558 1118
rect 1500 130 1512 1106
rect 1546 130 1558 1106
rect 1500 118 1558 130
rect -1558 -130 -1500 -118
rect -1558 -1106 -1546 -130
rect -1512 -1106 -1500 -130
rect -1558 -1118 -1500 -1106
rect 1500 -130 1558 -118
rect 1500 -1106 1512 -130
rect 1546 -1106 1558 -130
rect 1500 -1118 1558 -1106
rect -1558 -1366 -1500 -1354
rect -1558 -2342 -1546 -1366
rect -1512 -2342 -1500 -1366
rect -1558 -2354 -1500 -2342
rect 1500 -1366 1558 -1354
rect 1500 -2342 1512 -1366
rect 1546 -2342 1558 -1366
rect 1500 -2354 1558 -2342
rect -1558 -2602 -1500 -2590
rect -1558 -3578 -1546 -2602
rect -1512 -3578 -1500 -2602
rect -1558 -3590 -1500 -3578
rect 1500 -2602 1558 -2590
rect 1500 -3578 1512 -2602
rect 1546 -3578 1558 -2602
rect 1500 -3590 1558 -3578
rect -1558 -3838 -1500 -3826
rect -1558 -4814 -1546 -3838
rect -1512 -4814 -1500 -3838
rect -1558 -4826 -1500 -4814
rect 1500 -3838 1558 -3826
rect 1500 -4814 1512 -3838
rect 1546 -4814 1558 -3838
rect 1500 -4826 1558 -4814
rect -1558 -5074 -1500 -5062
rect -1558 -6050 -1546 -5074
rect -1512 -6050 -1500 -5074
rect -1558 -6062 -1500 -6050
rect 1500 -5074 1558 -5062
rect 1500 -6050 1512 -5074
rect 1546 -6050 1558 -5074
rect 1500 -6062 1558 -6050
rect -1558 -6310 -1500 -6298
rect -1558 -7286 -1546 -6310
rect -1512 -7286 -1500 -6310
rect -1558 -7298 -1500 -7286
rect 1500 -6310 1558 -6298
rect 1500 -7286 1512 -6310
rect 1546 -7286 1558 -6310
rect 1500 -7298 1558 -7286
rect -1558 -7546 -1500 -7534
rect -1558 -8522 -1546 -7546
rect -1512 -8522 -1500 -7546
rect -1558 -8534 -1500 -8522
rect 1500 -7546 1558 -7534
rect 1500 -8522 1512 -7546
rect 1546 -8522 1558 -7546
rect 1500 -8534 1558 -8522
rect -1558 -8782 -1500 -8770
rect -1558 -9758 -1546 -8782
rect -1512 -9758 -1500 -8782
rect -1558 -9770 -1500 -9758
rect 1500 -8782 1558 -8770
rect 1500 -9758 1512 -8782
rect 1546 -9758 1558 -8782
rect 1500 -9770 1558 -9758
rect -1558 -10018 -1500 -10006
rect -1558 -10994 -1546 -10018
rect -1512 -10994 -1500 -10018
rect -1558 -11006 -1500 -10994
rect 1500 -10018 1558 -10006
rect 1500 -10994 1512 -10018
rect 1546 -10994 1558 -10018
rect 1500 -11006 1558 -10994
rect -1558 -11254 -1500 -11242
rect -1558 -12230 -1546 -11254
rect -1512 -12230 -1500 -11254
rect -1558 -12242 -1500 -12230
rect 1500 -11254 1558 -11242
rect 1500 -12230 1512 -11254
rect 1546 -12230 1558 -11254
rect 1500 -12242 1558 -12230
rect -1558 -12490 -1500 -12478
rect -1558 -13466 -1546 -12490
rect -1512 -13466 -1500 -12490
rect -1558 -13478 -1500 -13466
rect 1500 -12490 1558 -12478
rect 1500 -13466 1512 -12490
rect 1546 -13466 1558 -12490
rect 1500 -13478 1558 -13466
rect -1558 -13726 -1500 -13714
rect -1558 -14702 -1546 -13726
rect -1512 -14702 -1500 -13726
rect -1558 -14714 -1500 -14702
rect 1500 -13726 1558 -13714
rect 1500 -14702 1512 -13726
rect 1546 -14702 1558 -13726
rect 1500 -14714 1558 -14702
rect -1558 -14962 -1500 -14950
rect -1558 -15938 -1546 -14962
rect -1512 -15938 -1500 -14962
rect -1558 -15950 -1500 -15938
rect 1500 -14962 1558 -14950
rect 1500 -15938 1512 -14962
rect 1546 -15938 1558 -14962
rect 1500 -15950 1558 -15938
rect -1558 -16198 -1500 -16186
rect -1558 -17174 -1546 -16198
rect -1512 -17174 -1500 -16198
rect -1558 -17186 -1500 -17174
rect 1500 -16198 1558 -16186
rect 1500 -17174 1512 -16198
rect 1546 -17174 1558 -16198
rect 1500 -17186 1558 -17174
rect -1558 -17434 -1500 -17422
rect -1558 -18410 -1546 -17434
rect -1512 -18410 -1500 -17434
rect -1558 -18422 -1500 -18410
rect 1500 -17434 1558 -17422
rect 1500 -18410 1512 -17434
rect 1546 -18410 1558 -17434
rect 1500 -18422 1558 -18410
rect -1558 -18670 -1500 -18658
rect -1558 -19646 -1546 -18670
rect -1512 -19646 -1500 -18670
rect -1558 -19658 -1500 -19646
rect 1500 -18670 1558 -18658
rect 1500 -19646 1512 -18670
rect 1546 -19646 1558 -18670
rect 1500 -19658 1558 -19646
rect -1558 -19906 -1500 -19894
rect -1558 -20882 -1546 -19906
rect -1512 -20882 -1500 -19906
rect -1558 -20894 -1500 -20882
rect 1500 -19906 1558 -19894
rect 1500 -20882 1512 -19906
rect 1546 -20882 1558 -19906
rect 1500 -20894 1558 -20882
rect -1558 -21142 -1500 -21130
rect -1558 -22118 -1546 -21142
rect -1512 -22118 -1500 -21142
rect -1558 -22130 -1500 -22118
rect 1500 -21142 1558 -21130
rect 1500 -22118 1512 -21142
rect 1546 -22118 1558 -21142
rect 1500 -22130 1558 -22118
rect -1558 -22378 -1500 -22366
rect -1558 -23354 -1546 -22378
rect -1512 -23354 -1500 -22378
rect -1558 -23366 -1500 -23354
rect 1500 -22378 1558 -22366
rect 1500 -23354 1512 -22378
rect 1546 -23354 1558 -22378
rect 1500 -23366 1558 -23354
rect -1558 -23614 -1500 -23602
rect -1558 -24590 -1546 -23614
rect -1512 -24590 -1500 -23614
rect -1558 -24602 -1500 -24590
rect 1500 -23614 1558 -23602
rect 1500 -24590 1512 -23614
rect 1546 -24590 1558 -23614
rect 1500 -24602 1558 -24590
rect -1558 -24850 -1500 -24838
rect -1558 -25826 -1546 -24850
rect -1512 -25826 -1500 -24850
rect -1558 -25838 -1500 -25826
rect 1500 -24850 1558 -24838
rect 1500 -25826 1512 -24850
rect 1546 -25826 1558 -24850
rect 1500 -25838 1558 -25826
rect -1558 -26086 -1500 -26074
rect -1558 -27062 -1546 -26086
rect -1512 -27062 -1500 -26086
rect -1558 -27074 -1500 -27062
rect 1500 -26086 1558 -26074
rect 1500 -27062 1512 -26086
rect 1546 -27062 1558 -26086
rect 1500 -27074 1558 -27062
rect -1558 -27322 -1500 -27310
rect -1558 -28298 -1546 -27322
rect -1512 -28298 -1500 -27322
rect -1558 -28310 -1500 -28298
rect 1500 -27322 1558 -27310
rect 1500 -28298 1512 -27322
rect 1546 -28298 1558 -27322
rect 1500 -28310 1558 -28298
rect -1558 -28558 -1500 -28546
rect -1558 -29534 -1546 -28558
rect -1512 -29534 -1500 -28558
rect -1558 -29546 -1500 -29534
rect 1500 -28558 1558 -28546
rect 1500 -29534 1512 -28558
rect 1546 -29534 1558 -28558
rect 1500 -29546 1558 -29534
rect -1558 -29794 -1500 -29782
rect -1558 -30770 -1546 -29794
rect -1512 -30770 -1500 -29794
rect -1558 -30782 -1500 -30770
rect 1500 -29794 1558 -29782
rect 1500 -30770 1512 -29794
rect 1546 -30770 1558 -29794
rect 1500 -30782 1558 -30770
rect -1558 -31030 -1500 -31018
rect -1558 -32006 -1546 -31030
rect -1512 -32006 -1500 -31030
rect -1558 -32018 -1500 -32006
rect 1500 -31030 1558 -31018
rect 1500 -32006 1512 -31030
rect 1546 -32006 1558 -31030
rect 1500 -32018 1558 -32006
rect -1558 -32266 -1500 -32254
rect -1558 -33242 -1546 -32266
rect -1512 -33242 -1500 -32266
rect -1558 -33254 -1500 -33242
rect 1500 -32266 1558 -32254
rect 1500 -33242 1512 -32266
rect 1546 -33242 1558 -32266
rect 1500 -33254 1558 -33242
rect -1558 -33502 -1500 -33490
rect -1558 -34478 -1546 -33502
rect -1512 -34478 -1500 -33502
rect -1558 -34490 -1500 -34478
rect 1500 -33502 1558 -33490
rect 1500 -34478 1512 -33502
rect 1546 -34478 1558 -33502
rect 1500 -34490 1558 -34478
rect -1558 -34738 -1500 -34726
rect -1558 -35714 -1546 -34738
rect -1512 -35714 -1500 -34738
rect -1558 -35726 -1500 -35714
rect 1500 -34738 1558 -34726
rect 1500 -35714 1512 -34738
rect 1546 -35714 1558 -34738
rect 1500 -35726 1558 -35714
rect -1558 -35974 -1500 -35962
rect -1558 -36950 -1546 -35974
rect -1512 -36950 -1500 -35974
rect -1558 -36962 -1500 -36950
rect 1500 -35974 1558 -35962
rect 1500 -36950 1512 -35974
rect 1546 -36950 1558 -35974
rect 1500 -36962 1558 -36950
rect -1558 -37210 -1500 -37198
rect -1558 -38186 -1546 -37210
rect -1512 -38186 -1500 -37210
rect -1558 -38198 -1500 -38186
rect 1500 -37210 1558 -37198
rect 1500 -38186 1512 -37210
rect 1546 -38186 1558 -37210
rect 1500 -38198 1558 -38186
rect -1558 -38446 -1500 -38434
rect -1558 -39422 -1546 -38446
rect -1512 -39422 -1500 -38446
rect -1558 -39434 -1500 -39422
rect 1500 -38446 1558 -38434
rect 1500 -39422 1512 -38446
rect 1546 -39422 1558 -38446
rect 1500 -39434 1558 -39422
rect -1558 -39682 -1500 -39670
rect -1558 -40658 -1546 -39682
rect -1512 -40658 -1500 -39682
rect -1558 -40670 -1500 -40658
rect 1500 -39682 1558 -39670
rect 1500 -40658 1512 -39682
rect 1546 -40658 1558 -39682
rect 1500 -40670 1558 -40658
rect -1558 -40918 -1500 -40906
rect -1558 -41894 -1546 -40918
rect -1512 -41894 -1500 -40918
rect -1558 -41906 -1500 -41894
rect 1500 -40918 1558 -40906
rect 1500 -41894 1512 -40918
rect 1546 -41894 1558 -40918
rect 1500 -41906 1558 -41894
rect -1558 -42154 -1500 -42142
rect -1558 -43130 -1546 -42154
rect -1512 -43130 -1500 -42154
rect -1558 -43142 -1500 -43130
rect 1500 -42154 1558 -42142
rect 1500 -43130 1512 -42154
rect 1546 -43130 1558 -42154
rect 1500 -43142 1558 -43130
rect -1558 -43390 -1500 -43378
rect -1558 -44366 -1546 -43390
rect -1512 -44366 -1500 -43390
rect -1558 -44378 -1500 -44366
rect 1500 -43390 1558 -43378
rect 1500 -44366 1512 -43390
rect 1546 -44366 1558 -43390
rect 1500 -44378 1558 -44366
rect -1558 -44626 -1500 -44614
rect -1558 -45602 -1546 -44626
rect -1512 -45602 -1500 -44626
rect -1558 -45614 -1500 -45602
rect 1500 -44626 1558 -44614
rect 1500 -45602 1512 -44626
rect 1546 -45602 1558 -44626
rect 1500 -45614 1558 -45602
rect -1558 -45862 -1500 -45850
rect -1558 -46838 -1546 -45862
rect -1512 -46838 -1500 -45862
rect -1558 -46850 -1500 -46838
rect 1500 -45862 1558 -45850
rect 1500 -46838 1512 -45862
rect 1546 -46838 1558 -45862
rect 1500 -46850 1558 -46838
rect -1558 -47098 -1500 -47086
rect -1558 -48074 -1546 -47098
rect -1512 -48074 -1500 -47098
rect -1558 -48086 -1500 -48074
rect 1500 -47098 1558 -47086
rect 1500 -48074 1512 -47098
rect 1546 -48074 1558 -47098
rect 1500 -48086 1558 -48074
rect -1558 -48334 -1500 -48322
rect -1558 -49310 -1546 -48334
rect -1512 -49310 -1500 -48334
rect -1558 -49322 -1500 -49310
rect 1500 -48334 1558 -48322
rect 1500 -49310 1512 -48334
rect 1546 -49310 1558 -48334
rect 1500 -49322 1558 -49310
rect -1558 -49570 -1500 -49558
rect -1558 -50546 -1546 -49570
rect -1512 -50546 -1500 -49570
rect -1558 -50558 -1500 -50546
rect 1500 -49570 1558 -49558
rect 1500 -50546 1512 -49570
rect 1546 -50546 1558 -49570
rect 1500 -50558 1558 -50546
rect -1558 -50806 -1500 -50794
rect -1558 -51782 -1546 -50806
rect -1512 -51782 -1500 -50806
rect -1558 -51794 -1500 -51782
rect 1500 -50806 1558 -50794
rect 1500 -51782 1512 -50806
rect 1546 -51782 1558 -50806
rect 1500 -51794 1558 -51782
rect -1558 -52042 -1500 -52030
rect -1558 -53018 -1546 -52042
rect -1512 -53018 -1500 -52042
rect -1558 -53030 -1500 -53018
rect 1500 -52042 1558 -52030
rect 1500 -53018 1512 -52042
rect 1546 -53018 1558 -52042
rect 1500 -53030 1558 -53018
rect -1558 -53278 -1500 -53266
rect -1558 -54254 -1546 -53278
rect -1512 -54254 -1500 -53278
rect -1558 -54266 -1500 -54254
rect 1500 -53278 1558 -53266
rect 1500 -54254 1512 -53278
rect 1546 -54254 1558 -53278
rect 1500 -54266 1558 -54254
rect -1558 -54514 -1500 -54502
rect -1558 -55490 -1546 -54514
rect -1512 -55490 -1500 -54514
rect -1558 -55502 -1500 -55490
rect 1500 -54514 1558 -54502
rect 1500 -55490 1512 -54514
rect 1546 -55490 1558 -54514
rect 1500 -55502 1558 -55490
rect -1558 -55750 -1500 -55738
rect -1558 -56726 -1546 -55750
rect -1512 -56726 -1500 -55750
rect -1558 -56738 -1500 -56726
rect 1500 -55750 1558 -55738
rect 1500 -56726 1512 -55750
rect 1546 -56726 1558 -55750
rect 1500 -56738 1558 -56726
rect -1558 -56986 -1500 -56974
rect -1558 -57962 -1546 -56986
rect -1512 -57962 -1500 -56986
rect -1558 -57974 -1500 -57962
rect 1500 -56986 1558 -56974
rect 1500 -57962 1512 -56986
rect 1546 -57962 1558 -56986
rect 1500 -57974 1558 -57962
rect -1558 -58222 -1500 -58210
rect -1558 -59198 -1546 -58222
rect -1512 -59198 -1500 -58222
rect -1558 -59210 -1500 -59198
rect 1500 -58222 1558 -58210
rect 1500 -59198 1512 -58222
rect 1546 -59198 1558 -58222
rect 1500 -59210 1558 -59198
rect -1558 -59458 -1500 -59446
rect -1558 -60434 -1546 -59458
rect -1512 -60434 -1500 -59458
rect -1558 -60446 -1500 -60434
rect 1500 -59458 1558 -59446
rect 1500 -60434 1512 -59458
rect 1546 -60434 1558 -59458
rect 1500 -60446 1558 -60434
rect -1558 -60694 -1500 -60682
rect -1558 -61670 -1546 -60694
rect -1512 -61670 -1500 -60694
rect -1558 -61682 -1500 -61670
rect 1500 -60694 1558 -60682
rect 1500 -61670 1512 -60694
rect 1546 -61670 1558 -60694
rect 1500 -61682 1558 -61670
rect -1558 -61930 -1500 -61918
rect -1558 -62906 -1546 -61930
rect -1512 -62906 -1500 -61930
rect -1558 -62918 -1500 -62906
rect 1500 -61930 1558 -61918
rect 1500 -62906 1512 -61930
rect 1546 -62906 1558 -61930
rect 1500 -62918 1558 -62906
<< pdiffc >>
rect -1546 61930 -1512 62906
rect 1512 61930 1546 62906
rect -1546 60694 -1512 61670
rect 1512 60694 1546 61670
rect -1546 59458 -1512 60434
rect 1512 59458 1546 60434
rect -1546 58222 -1512 59198
rect 1512 58222 1546 59198
rect -1546 56986 -1512 57962
rect 1512 56986 1546 57962
rect -1546 55750 -1512 56726
rect 1512 55750 1546 56726
rect -1546 54514 -1512 55490
rect 1512 54514 1546 55490
rect -1546 53278 -1512 54254
rect 1512 53278 1546 54254
rect -1546 52042 -1512 53018
rect 1512 52042 1546 53018
rect -1546 50806 -1512 51782
rect 1512 50806 1546 51782
rect -1546 49570 -1512 50546
rect 1512 49570 1546 50546
rect -1546 48334 -1512 49310
rect 1512 48334 1546 49310
rect -1546 47098 -1512 48074
rect 1512 47098 1546 48074
rect -1546 45862 -1512 46838
rect 1512 45862 1546 46838
rect -1546 44626 -1512 45602
rect 1512 44626 1546 45602
rect -1546 43390 -1512 44366
rect 1512 43390 1546 44366
rect -1546 42154 -1512 43130
rect 1512 42154 1546 43130
rect -1546 40918 -1512 41894
rect 1512 40918 1546 41894
rect -1546 39682 -1512 40658
rect 1512 39682 1546 40658
rect -1546 38446 -1512 39422
rect 1512 38446 1546 39422
rect -1546 37210 -1512 38186
rect 1512 37210 1546 38186
rect -1546 35974 -1512 36950
rect 1512 35974 1546 36950
rect -1546 34738 -1512 35714
rect 1512 34738 1546 35714
rect -1546 33502 -1512 34478
rect 1512 33502 1546 34478
rect -1546 32266 -1512 33242
rect 1512 32266 1546 33242
rect -1546 31030 -1512 32006
rect 1512 31030 1546 32006
rect -1546 29794 -1512 30770
rect 1512 29794 1546 30770
rect -1546 28558 -1512 29534
rect 1512 28558 1546 29534
rect -1546 27322 -1512 28298
rect 1512 27322 1546 28298
rect -1546 26086 -1512 27062
rect 1512 26086 1546 27062
rect -1546 24850 -1512 25826
rect 1512 24850 1546 25826
rect -1546 23614 -1512 24590
rect 1512 23614 1546 24590
rect -1546 22378 -1512 23354
rect 1512 22378 1546 23354
rect -1546 21142 -1512 22118
rect 1512 21142 1546 22118
rect -1546 19906 -1512 20882
rect 1512 19906 1546 20882
rect -1546 18670 -1512 19646
rect 1512 18670 1546 19646
rect -1546 17434 -1512 18410
rect 1512 17434 1546 18410
rect -1546 16198 -1512 17174
rect 1512 16198 1546 17174
rect -1546 14962 -1512 15938
rect 1512 14962 1546 15938
rect -1546 13726 -1512 14702
rect 1512 13726 1546 14702
rect -1546 12490 -1512 13466
rect 1512 12490 1546 13466
rect -1546 11254 -1512 12230
rect 1512 11254 1546 12230
rect -1546 10018 -1512 10994
rect 1512 10018 1546 10994
rect -1546 8782 -1512 9758
rect 1512 8782 1546 9758
rect -1546 7546 -1512 8522
rect 1512 7546 1546 8522
rect -1546 6310 -1512 7286
rect 1512 6310 1546 7286
rect -1546 5074 -1512 6050
rect 1512 5074 1546 6050
rect -1546 3838 -1512 4814
rect 1512 3838 1546 4814
rect -1546 2602 -1512 3578
rect 1512 2602 1546 3578
rect -1546 1366 -1512 2342
rect 1512 1366 1546 2342
rect -1546 130 -1512 1106
rect 1512 130 1546 1106
rect -1546 -1106 -1512 -130
rect 1512 -1106 1546 -130
rect -1546 -2342 -1512 -1366
rect 1512 -2342 1546 -1366
rect -1546 -3578 -1512 -2602
rect 1512 -3578 1546 -2602
rect -1546 -4814 -1512 -3838
rect 1512 -4814 1546 -3838
rect -1546 -6050 -1512 -5074
rect 1512 -6050 1546 -5074
rect -1546 -7286 -1512 -6310
rect 1512 -7286 1546 -6310
rect -1546 -8522 -1512 -7546
rect 1512 -8522 1546 -7546
rect -1546 -9758 -1512 -8782
rect 1512 -9758 1546 -8782
rect -1546 -10994 -1512 -10018
rect 1512 -10994 1546 -10018
rect -1546 -12230 -1512 -11254
rect 1512 -12230 1546 -11254
rect -1546 -13466 -1512 -12490
rect 1512 -13466 1546 -12490
rect -1546 -14702 -1512 -13726
rect 1512 -14702 1546 -13726
rect -1546 -15938 -1512 -14962
rect 1512 -15938 1546 -14962
rect -1546 -17174 -1512 -16198
rect 1512 -17174 1546 -16198
rect -1546 -18410 -1512 -17434
rect 1512 -18410 1546 -17434
rect -1546 -19646 -1512 -18670
rect 1512 -19646 1546 -18670
rect -1546 -20882 -1512 -19906
rect 1512 -20882 1546 -19906
rect -1546 -22118 -1512 -21142
rect 1512 -22118 1546 -21142
rect -1546 -23354 -1512 -22378
rect 1512 -23354 1546 -22378
rect -1546 -24590 -1512 -23614
rect 1512 -24590 1546 -23614
rect -1546 -25826 -1512 -24850
rect 1512 -25826 1546 -24850
rect -1546 -27062 -1512 -26086
rect 1512 -27062 1546 -26086
rect -1546 -28298 -1512 -27322
rect 1512 -28298 1546 -27322
rect -1546 -29534 -1512 -28558
rect 1512 -29534 1546 -28558
rect -1546 -30770 -1512 -29794
rect 1512 -30770 1546 -29794
rect -1546 -32006 -1512 -31030
rect 1512 -32006 1546 -31030
rect -1546 -33242 -1512 -32266
rect 1512 -33242 1546 -32266
rect -1546 -34478 -1512 -33502
rect 1512 -34478 1546 -33502
rect -1546 -35714 -1512 -34738
rect 1512 -35714 1546 -34738
rect -1546 -36950 -1512 -35974
rect 1512 -36950 1546 -35974
rect -1546 -38186 -1512 -37210
rect 1512 -38186 1546 -37210
rect -1546 -39422 -1512 -38446
rect 1512 -39422 1546 -38446
rect -1546 -40658 -1512 -39682
rect 1512 -40658 1546 -39682
rect -1546 -41894 -1512 -40918
rect 1512 -41894 1546 -40918
rect -1546 -43130 -1512 -42154
rect 1512 -43130 1546 -42154
rect -1546 -44366 -1512 -43390
rect 1512 -44366 1546 -43390
rect -1546 -45602 -1512 -44626
rect 1512 -45602 1546 -44626
rect -1546 -46838 -1512 -45862
rect 1512 -46838 1546 -45862
rect -1546 -48074 -1512 -47098
rect 1512 -48074 1546 -47098
rect -1546 -49310 -1512 -48334
rect 1512 -49310 1546 -48334
rect -1546 -50546 -1512 -49570
rect 1512 -50546 1546 -49570
rect -1546 -51782 -1512 -50806
rect 1512 -51782 1546 -50806
rect -1546 -53018 -1512 -52042
rect 1512 -53018 1546 -52042
rect -1546 -54254 -1512 -53278
rect 1512 -54254 1546 -53278
rect -1546 -55490 -1512 -54514
rect 1512 -55490 1546 -54514
rect -1546 -56726 -1512 -55750
rect 1512 -56726 1546 -55750
rect -1546 -57962 -1512 -56986
rect 1512 -57962 1546 -56986
rect -1546 -59198 -1512 -58222
rect 1512 -59198 1546 -58222
rect -1546 -60434 -1512 -59458
rect 1512 -60434 1546 -59458
rect -1546 -61670 -1512 -60694
rect 1512 -61670 1546 -60694
rect -1546 -62906 -1512 -61930
rect 1512 -62906 1546 -61930
<< poly >>
rect -1500 62999 1500 63015
rect -1500 62965 -1484 62999
rect 1484 62965 1500 62999
rect -1500 62918 1500 62965
rect -1500 61871 1500 61918
rect -1500 61837 -1484 61871
rect 1484 61837 1500 61871
rect -1500 61821 1500 61837
rect -1500 61763 1500 61779
rect -1500 61729 -1484 61763
rect 1484 61729 1500 61763
rect -1500 61682 1500 61729
rect -1500 60635 1500 60682
rect -1500 60601 -1484 60635
rect 1484 60601 1500 60635
rect -1500 60585 1500 60601
rect -1500 60527 1500 60543
rect -1500 60493 -1484 60527
rect 1484 60493 1500 60527
rect -1500 60446 1500 60493
rect -1500 59399 1500 59446
rect -1500 59365 -1484 59399
rect 1484 59365 1500 59399
rect -1500 59349 1500 59365
rect -1500 59291 1500 59307
rect -1500 59257 -1484 59291
rect 1484 59257 1500 59291
rect -1500 59210 1500 59257
rect -1500 58163 1500 58210
rect -1500 58129 -1484 58163
rect 1484 58129 1500 58163
rect -1500 58113 1500 58129
rect -1500 58055 1500 58071
rect -1500 58021 -1484 58055
rect 1484 58021 1500 58055
rect -1500 57974 1500 58021
rect -1500 56927 1500 56974
rect -1500 56893 -1484 56927
rect 1484 56893 1500 56927
rect -1500 56877 1500 56893
rect -1500 56819 1500 56835
rect -1500 56785 -1484 56819
rect 1484 56785 1500 56819
rect -1500 56738 1500 56785
rect -1500 55691 1500 55738
rect -1500 55657 -1484 55691
rect 1484 55657 1500 55691
rect -1500 55641 1500 55657
rect -1500 55583 1500 55599
rect -1500 55549 -1484 55583
rect 1484 55549 1500 55583
rect -1500 55502 1500 55549
rect -1500 54455 1500 54502
rect -1500 54421 -1484 54455
rect 1484 54421 1500 54455
rect -1500 54405 1500 54421
rect -1500 54347 1500 54363
rect -1500 54313 -1484 54347
rect 1484 54313 1500 54347
rect -1500 54266 1500 54313
rect -1500 53219 1500 53266
rect -1500 53185 -1484 53219
rect 1484 53185 1500 53219
rect -1500 53169 1500 53185
rect -1500 53111 1500 53127
rect -1500 53077 -1484 53111
rect 1484 53077 1500 53111
rect -1500 53030 1500 53077
rect -1500 51983 1500 52030
rect -1500 51949 -1484 51983
rect 1484 51949 1500 51983
rect -1500 51933 1500 51949
rect -1500 51875 1500 51891
rect -1500 51841 -1484 51875
rect 1484 51841 1500 51875
rect -1500 51794 1500 51841
rect -1500 50747 1500 50794
rect -1500 50713 -1484 50747
rect 1484 50713 1500 50747
rect -1500 50697 1500 50713
rect -1500 50639 1500 50655
rect -1500 50605 -1484 50639
rect 1484 50605 1500 50639
rect -1500 50558 1500 50605
rect -1500 49511 1500 49558
rect -1500 49477 -1484 49511
rect 1484 49477 1500 49511
rect -1500 49461 1500 49477
rect -1500 49403 1500 49419
rect -1500 49369 -1484 49403
rect 1484 49369 1500 49403
rect -1500 49322 1500 49369
rect -1500 48275 1500 48322
rect -1500 48241 -1484 48275
rect 1484 48241 1500 48275
rect -1500 48225 1500 48241
rect -1500 48167 1500 48183
rect -1500 48133 -1484 48167
rect 1484 48133 1500 48167
rect -1500 48086 1500 48133
rect -1500 47039 1500 47086
rect -1500 47005 -1484 47039
rect 1484 47005 1500 47039
rect -1500 46989 1500 47005
rect -1500 46931 1500 46947
rect -1500 46897 -1484 46931
rect 1484 46897 1500 46931
rect -1500 46850 1500 46897
rect -1500 45803 1500 45850
rect -1500 45769 -1484 45803
rect 1484 45769 1500 45803
rect -1500 45753 1500 45769
rect -1500 45695 1500 45711
rect -1500 45661 -1484 45695
rect 1484 45661 1500 45695
rect -1500 45614 1500 45661
rect -1500 44567 1500 44614
rect -1500 44533 -1484 44567
rect 1484 44533 1500 44567
rect -1500 44517 1500 44533
rect -1500 44459 1500 44475
rect -1500 44425 -1484 44459
rect 1484 44425 1500 44459
rect -1500 44378 1500 44425
rect -1500 43331 1500 43378
rect -1500 43297 -1484 43331
rect 1484 43297 1500 43331
rect -1500 43281 1500 43297
rect -1500 43223 1500 43239
rect -1500 43189 -1484 43223
rect 1484 43189 1500 43223
rect -1500 43142 1500 43189
rect -1500 42095 1500 42142
rect -1500 42061 -1484 42095
rect 1484 42061 1500 42095
rect -1500 42045 1500 42061
rect -1500 41987 1500 42003
rect -1500 41953 -1484 41987
rect 1484 41953 1500 41987
rect -1500 41906 1500 41953
rect -1500 40859 1500 40906
rect -1500 40825 -1484 40859
rect 1484 40825 1500 40859
rect -1500 40809 1500 40825
rect -1500 40751 1500 40767
rect -1500 40717 -1484 40751
rect 1484 40717 1500 40751
rect -1500 40670 1500 40717
rect -1500 39623 1500 39670
rect -1500 39589 -1484 39623
rect 1484 39589 1500 39623
rect -1500 39573 1500 39589
rect -1500 39515 1500 39531
rect -1500 39481 -1484 39515
rect 1484 39481 1500 39515
rect -1500 39434 1500 39481
rect -1500 38387 1500 38434
rect -1500 38353 -1484 38387
rect 1484 38353 1500 38387
rect -1500 38337 1500 38353
rect -1500 38279 1500 38295
rect -1500 38245 -1484 38279
rect 1484 38245 1500 38279
rect -1500 38198 1500 38245
rect -1500 37151 1500 37198
rect -1500 37117 -1484 37151
rect 1484 37117 1500 37151
rect -1500 37101 1500 37117
rect -1500 37043 1500 37059
rect -1500 37009 -1484 37043
rect 1484 37009 1500 37043
rect -1500 36962 1500 37009
rect -1500 35915 1500 35962
rect -1500 35881 -1484 35915
rect 1484 35881 1500 35915
rect -1500 35865 1500 35881
rect -1500 35807 1500 35823
rect -1500 35773 -1484 35807
rect 1484 35773 1500 35807
rect -1500 35726 1500 35773
rect -1500 34679 1500 34726
rect -1500 34645 -1484 34679
rect 1484 34645 1500 34679
rect -1500 34629 1500 34645
rect -1500 34571 1500 34587
rect -1500 34537 -1484 34571
rect 1484 34537 1500 34571
rect -1500 34490 1500 34537
rect -1500 33443 1500 33490
rect -1500 33409 -1484 33443
rect 1484 33409 1500 33443
rect -1500 33393 1500 33409
rect -1500 33335 1500 33351
rect -1500 33301 -1484 33335
rect 1484 33301 1500 33335
rect -1500 33254 1500 33301
rect -1500 32207 1500 32254
rect -1500 32173 -1484 32207
rect 1484 32173 1500 32207
rect -1500 32157 1500 32173
rect -1500 32099 1500 32115
rect -1500 32065 -1484 32099
rect 1484 32065 1500 32099
rect -1500 32018 1500 32065
rect -1500 30971 1500 31018
rect -1500 30937 -1484 30971
rect 1484 30937 1500 30971
rect -1500 30921 1500 30937
rect -1500 30863 1500 30879
rect -1500 30829 -1484 30863
rect 1484 30829 1500 30863
rect -1500 30782 1500 30829
rect -1500 29735 1500 29782
rect -1500 29701 -1484 29735
rect 1484 29701 1500 29735
rect -1500 29685 1500 29701
rect -1500 29627 1500 29643
rect -1500 29593 -1484 29627
rect 1484 29593 1500 29627
rect -1500 29546 1500 29593
rect -1500 28499 1500 28546
rect -1500 28465 -1484 28499
rect 1484 28465 1500 28499
rect -1500 28449 1500 28465
rect -1500 28391 1500 28407
rect -1500 28357 -1484 28391
rect 1484 28357 1500 28391
rect -1500 28310 1500 28357
rect -1500 27263 1500 27310
rect -1500 27229 -1484 27263
rect 1484 27229 1500 27263
rect -1500 27213 1500 27229
rect -1500 27155 1500 27171
rect -1500 27121 -1484 27155
rect 1484 27121 1500 27155
rect -1500 27074 1500 27121
rect -1500 26027 1500 26074
rect -1500 25993 -1484 26027
rect 1484 25993 1500 26027
rect -1500 25977 1500 25993
rect -1500 25919 1500 25935
rect -1500 25885 -1484 25919
rect 1484 25885 1500 25919
rect -1500 25838 1500 25885
rect -1500 24791 1500 24838
rect -1500 24757 -1484 24791
rect 1484 24757 1500 24791
rect -1500 24741 1500 24757
rect -1500 24683 1500 24699
rect -1500 24649 -1484 24683
rect 1484 24649 1500 24683
rect -1500 24602 1500 24649
rect -1500 23555 1500 23602
rect -1500 23521 -1484 23555
rect 1484 23521 1500 23555
rect -1500 23505 1500 23521
rect -1500 23447 1500 23463
rect -1500 23413 -1484 23447
rect 1484 23413 1500 23447
rect -1500 23366 1500 23413
rect -1500 22319 1500 22366
rect -1500 22285 -1484 22319
rect 1484 22285 1500 22319
rect -1500 22269 1500 22285
rect -1500 22211 1500 22227
rect -1500 22177 -1484 22211
rect 1484 22177 1500 22211
rect -1500 22130 1500 22177
rect -1500 21083 1500 21130
rect -1500 21049 -1484 21083
rect 1484 21049 1500 21083
rect -1500 21033 1500 21049
rect -1500 20975 1500 20991
rect -1500 20941 -1484 20975
rect 1484 20941 1500 20975
rect -1500 20894 1500 20941
rect -1500 19847 1500 19894
rect -1500 19813 -1484 19847
rect 1484 19813 1500 19847
rect -1500 19797 1500 19813
rect -1500 19739 1500 19755
rect -1500 19705 -1484 19739
rect 1484 19705 1500 19739
rect -1500 19658 1500 19705
rect -1500 18611 1500 18658
rect -1500 18577 -1484 18611
rect 1484 18577 1500 18611
rect -1500 18561 1500 18577
rect -1500 18503 1500 18519
rect -1500 18469 -1484 18503
rect 1484 18469 1500 18503
rect -1500 18422 1500 18469
rect -1500 17375 1500 17422
rect -1500 17341 -1484 17375
rect 1484 17341 1500 17375
rect -1500 17325 1500 17341
rect -1500 17267 1500 17283
rect -1500 17233 -1484 17267
rect 1484 17233 1500 17267
rect -1500 17186 1500 17233
rect -1500 16139 1500 16186
rect -1500 16105 -1484 16139
rect 1484 16105 1500 16139
rect -1500 16089 1500 16105
rect -1500 16031 1500 16047
rect -1500 15997 -1484 16031
rect 1484 15997 1500 16031
rect -1500 15950 1500 15997
rect -1500 14903 1500 14950
rect -1500 14869 -1484 14903
rect 1484 14869 1500 14903
rect -1500 14853 1500 14869
rect -1500 14795 1500 14811
rect -1500 14761 -1484 14795
rect 1484 14761 1500 14795
rect -1500 14714 1500 14761
rect -1500 13667 1500 13714
rect -1500 13633 -1484 13667
rect 1484 13633 1500 13667
rect -1500 13617 1500 13633
rect -1500 13559 1500 13575
rect -1500 13525 -1484 13559
rect 1484 13525 1500 13559
rect -1500 13478 1500 13525
rect -1500 12431 1500 12478
rect -1500 12397 -1484 12431
rect 1484 12397 1500 12431
rect -1500 12381 1500 12397
rect -1500 12323 1500 12339
rect -1500 12289 -1484 12323
rect 1484 12289 1500 12323
rect -1500 12242 1500 12289
rect -1500 11195 1500 11242
rect -1500 11161 -1484 11195
rect 1484 11161 1500 11195
rect -1500 11145 1500 11161
rect -1500 11087 1500 11103
rect -1500 11053 -1484 11087
rect 1484 11053 1500 11087
rect -1500 11006 1500 11053
rect -1500 9959 1500 10006
rect -1500 9925 -1484 9959
rect 1484 9925 1500 9959
rect -1500 9909 1500 9925
rect -1500 9851 1500 9867
rect -1500 9817 -1484 9851
rect 1484 9817 1500 9851
rect -1500 9770 1500 9817
rect -1500 8723 1500 8770
rect -1500 8689 -1484 8723
rect 1484 8689 1500 8723
rect -1500 8673 1500 8689
rect -1500 8615 1500 8631
rect -1500 8581 -1484 8615
rect 1484 8581 1500 8615
rect -1500 8534 1500 8581
rect -1500 7487 1500 7534
rect -1500 7453 -1484 7487
rect 1484 7453 1500 7487
rect -1500 7437 1500 7453
rect -1500 7379 1500 7395
rect -1500 7345 -1484 7379
rect 1484 7345 1500 7379
rect -1500 7298 1500 7345
rect -1500 6251 1500 6298
rect -1500 6217 -1484 6251
rect 1484 6217 1500 6251
rect -1500 6201 1500 6217
rect -1500 6143 1500 6159
rect -1500 6109 -1484 6143
rect 1484 6109 1500 6143
rect -1500 6062 1500 6109
rect -1500 5015 1500 5062
rect -1500 4981 -1484 5015
rect 1484 4981 1500 5015
rect -1500 4965 1500 4981
rect -1500 4907 1500 4923
rect -1500 4873 -1484 4907
rect 1484 4873 1500 4907
rect -1500 4826 1500 4873
rect -1500 3779 1500 3826
rect -1500 3745 -1484 3779
rect 1484 3745 1500 3779
rect -1500 3729 1500 3745
rect -1500 3671 1500 3687
rect -1500 3637 -1484 3671
rect 1484 3637 1500 3671
rect -1500 3590 1500 3637
rect -1500 2543 1500 2590
rect -1500 2509 -1484 2543
rect 1484 2509 1500 2543
rect -1500 2493 1500 2509
rect -1500 2435 1500 2451
rect -1500 2401 -1484 2435
rect 1484 2401 1500 2435
rect -1500 2354 1500 2401
rect -1500 1307 1500 1354
rect -1500 1273 -1484 1307
rect 1484 1273 1500 1307
rect -1500 1257 1500 1273
rect -1500 1199 1500 1215
rect -1500 1165 -1484 1199
rect 1484 1165 1500 1199
rect -1500 1118 1500 1165
rect -1500 71 1500 118
rect -1500 37 -1484 71
rect 1484 37 1500 71
rect -1500 21 1500 37
rect -1500 -37 1500 -21
rect -1500 -71 -1484 -37
rect 1484 -71 1500 -37
rect -1500 -118 1500 -71
rect -1500 -1165 1500 -1118
rect -1500 -1199 -1484 -1165
rect 1484 -1199 1500 -1165
rect -1500 -1215 1500 -1199
rect -1500 -1273 1500 -1257
rect -1500 -1307 -1484 -1273
rect 1484 -1307 1500 -1273
rect -1500 -1354 1500 -1307
rect -1500 -2401 1500 -2354
rect -1500 -2435 -1484 -2401
rect 1484 -2435 1500 -2401
rect -1500 -2451 1500 -2435
rect -1500 -2509 1500 -2493
rect -1500 -2543 -1484 -2509
rect 1484 -2543 1500 -2509
rect -1500 -2590 1500 -2543
rect -1500 -3637 1500 -3590
rect -1500 -3671 -1484 -3637
rect 1484 -3671 1500 -3637
rect -1500 -3687 1500 -3671
rect -1500 -3745 1500 -3729
rect -1500 -3779 -1484 -3745
rect 1484 -3779 1500 -3745
rect -1500 -3826 1500 -3779
rect -1500 -4873 1500 -4826
rect -1500 -4907 -1484 -4873
rect 1484 -4907 1500 -4873
rect -1500 -4923 1500 -4907
rect -1500 -4981 1500 -4965
rect -1500 -5015 -1484 -4981
rect 1484 -5015 1500 -4981
rect -1500 -5062 1500 -5015
rect -1500 -6109 1500 -6062
rect -1500 -6143 -1484 -6109
rect 1484 -6143 1500 -6109
rect -1500 -6159 1500 -6143
rect -1500 -6217 1500 -6201
rect -1500 -6251 -1484 -6217
rect 1484 -6251 1500 -6217
rect -1500 -6298 1500 -6251
rect -1500 -7345 1500 -7298
rect -1500 -7379 -1484 -7345
rect 1484 -7379 1500 -7345
rect -1500 -7395 1500 -7379
rect -1500 -7453 1500 -7437
rect -1500 -7487 -1484 -7453
rect 1484 -7487 1500 -7453
rect -1500 -7534 1500 -7487
rect -1500 -8581 1500 -8534
rect -1500 -8615 -1484 -8581
rect 1484 -8615 1500 -8581
rect -1500 -8631 1500 -8615
rect -1500 -8689 1500 -8673
rect -1500 -8723 -1484 -8689
rect 1484 -8723 1500 -8689
rect -1500 -8770 1500 -8723
rect -1500 -9817 1500 -9770
rect -1500 -9851 -1484 -9817
rect 1484 -9851 1500 -9817
rect -1500 -9867 1500 -9851
rect -1500 -9925 1500 -9909
rect -1500 -9959 -1484 -9925
rect 1484 -9959 1500 -9925
rect -1500 -10006 1500 -9959
rect -1500 -11053 1500 -11006
rect -1500 -11087 -1484 -11053
rect 1484 -11087 1500 -11053
rect -1500 -11103 1500 -11087
rect -1500 -11161 1500 -11145
rect -1500 -11195 -1484 -11161
rect 1484 -11195 1500 -11161
rect -1500 -11242 1500 -11195
rect -1500 -12289 1500 -12242
rect -1500 -12323 -1484 -12289
rect 1484 -12323 1500 -12289
rect -1500 -12339 1500 -12323
rect -1500 -12397 1500 -12381
rect -1500 -12431 -1484 -12397
rect 1484 -12431 1500 -12397
rect -1500 -12478 1500 -12431
rect -1500 -13525 1500 -13478
rect -1500 -13559 -1484 -13525
rect 1484 -13559 1500 -13525
rect -1500 -13575 1500 -13559
rect -1500 -13633 1500 -13617
rect -1500 -13667 -1484 -13633
rect 1484 -13667 1500 -13633
rect -1500 -13714 1500 -13667
rect -1500 -14761 1500 -14714
rect -1500 -14795 -1484 -14761
rect 1484 -14795 1500 -14761
rect -1500 -14811 1500 -14795
rect -1500 -14869 1500 -14853
rect -1500 -14903 -1484 -14869
rect 1484 -14903 1500 -14869
rect -1500 -14950 1500 -14903
rect -1500 -15997 1500 -15950
rect -1500 -16031 -1484 -15997
rect 1484 -16031 1500 -15997
rect -1500 -16047 1500 -16031
rect -1500 -16105 1500 -16089
rect -1500 -16139 -1484 -16105
rect 1484 -16139 1500 -16105
rect -1500 -16186 1500 -16139
rect -1500 -17233 1500 -17186
rect -1500 -17267 -1484 -17233
rect 1484 -17267 1500 -17233
rect -1500 -17283 1500 -17267
rect -1500 -17341 1500 -17325
rect -1500 -17375 -1484 -17341
rect 1484 -17375 1500 -17341
rect -1500 -17422 1500 -17375
rect -1500 -18469 1500 -18422
rect -1500 -18503 -1484 -18469
rect 1484 -18503 1500 -18469
rect -1500 -18519 1500 -18503
rect -1500 -18577 1500 -18561
rect -1500 -18611 -1484 -18577
rect 1484 -18611 1500 -18577
rect -1500 -18658 1500 -18611
rect -1500 -19705 1500 -19658
rect -1500 -19739 -1484 -19705
rect 1484 -19739 1500 -19705
rect -1500 -19755 1500 -19739
rect -1500 -19813 1500 -19797
rect -1500 -19847 -1484 -19813
rect 1484 -19847 1500 -19813
rect -1500 -19894 1500 -19847
rect -1500 -20941 1500 -20894
rect -1500 -20975 -1484 -20941
rect 1484 -20975 1500 -20941
rect -1500 -20991 1500 -20975
rect -1500 -21049 1500 -21033
rect -1500 -21083 -1484 -21049
rect 1484 -21083 1500 -21049
rect -1500 -21130 1500 -21083
rect -1500 -22177 1500 -22130
rect -1500 -22211 -1484 -22177
rect 1484 -22211 1500 -22177
rect -1500 -22227 1500 -22211
rect -1500 -22285 1500 -22269
rect -1500 -22319 -1484 -22285
rect 1484 -22319 1500 -22285
rect -1500 -22366 1500 -22319
rect -1500 -23413 1500 -23366
rect -1500 -23447 -1484 -23413
rect 1484 -23447 1500 -23413
rect -1500 -23463 1500 -23447
rect -1500 -23521 1500 -23505
rect -1500 -23555 -1484 -23521
rect 1484 -23555 1500 -23521
rect -1500 -23602 1500 -23555
rect -1500 -24649 1500 -24602
rect -1500 -24683 -1484 -24649
rect 1484 -24683 1500 -24649
rect -1500 -24699 1500 -24683
rect -1500 -24757 1500 -24741
rect -1500 -24791 -1484 -24757
rect 1484 -24791 1500 -24757
rect -1500 -24838 1500 -24791
rect -1500 -25885 1500 -25838
rect -1500 -25919 -1484 -25885
rect 1484 -25919 1500 -25885
rect -1500 -25935 1500 -25919
rect -1500 -25993 1500 -25977
rect -1500 -26027 -1484 -25993
rect 1484 -26027 1500 -25993
rect -1500 -26074 1500 -26027
rect -1500 -27121 1500 -27074
rect -1500 -27155 -1484 -27121
rect 1484 -27155 1500 -27121
rect -1500 -27171 1500 -27155
rect -1500 -27229 1500 -27213
rect -1500 -27263 -1484 -27229
rect 1484 -27263 1500 -27229
rect -1500 -27310 1500 -27263
rect -1500 -28357 1500 -28310
rect -1500 -28391 -1484 -28357
rect 1484 -28391 1500 -28357
rect -1500 -28407 1500 -28391
rect -1500 -28465 1500 -28449
rect -1500 -28499 -1484 -28465
rect 1484 -28499 1500 -28465
rect -1500 -28546 1500 -28499
rect -1500 -29593 1500 -29546
rect -1500 -29627 -1484 -29593
rect 1484 -29627 1500 -29593
rect -1500 -29643 1500 -29627
rect -1500 -29701 1500 -29685
rect -1500 -29735 -1484 -29701
rect 1484 -29735 1500 -29701
rect -1500 -29782 1500 -29735
rect -1500 -30829 1500 -30782
rect -1500 -30863 -1484 -30829
rect 1484 -30863 1500 -30829
rect -1500 -30879 1500 -30863
rect -1500 -30937 1500 -30921
rect -1500 -30971 -1484 -30937
rect 1484 -30971 1500 -30937
rect -1500 -31018 1500 -30971
rect -1500 -32065 1500 -32018
rect -1500 -32099 -1484 -32065
rect 1484 -32099 1500 -32065
rect -1500 -32115 1500 -32099
rect -1500 -32173 1500 -32157
rect -1500 -32207 -1484 -32173
rect 1484 -32207 1500 -32173
rect -1500 -32254 1500 -32207
rect -1500 -33301 1500 -33254
rect -1500 -33335 -1484 -33301
rect 1484 -33335 1500 -33301
rect -1500 -33351 1500 -33335
rect -1500 -33409 1500 -33393
rect -1500 -33443 -1484 -33409
rect 1484 -33443 1500 -33409
rect -1500 -33490 1500 -33443
rect -1500 -34537 1500 -34490
rect -1500 -34571 -1484 -34537
rect 1484 -34571 1500 -34537
rect -1500 -34587 1500 -34571
rect -1500 -34645 1500 -34629
rect -1500 -34679 -1484 -34645
rect 1484 -34679 1500 -34645
rect -1500 -34726 1500 -34679
rect -1500 -35773 1500 -35726
rect -1500 -35807 -1484 -35773
rect 1484 -35807 1500 -35773
rect -1500 -35823 1500 -35807
rect -1500 -35881 1500 -35865
rect -1500 -35915 -1484 -35881
rect 1484 -35915 1500 -35881
rect -1500 -35962 1500 -35915
rect -1500 -37009 1500 -36962
rect -1500 -37043 -1484 -37009
rect 1484 -37043 1500 -37009
rect -1500 -37059 1500 -37043
rect -1500 -37117 1500 -37101
rect -1500 -37151 -1484 -37117
rect 1484 -37151 1500 -37117
rect -1500 -37198 1500 -37151
rect -1500 -38245 1500 -38198
rect -1500 -38279 -1484 -38245
rect 1484 -38279 1500 -38245
rect -1500 -38295 1500 -38279
rect -1500 -38353 1500 -38337
rect -1500 -38387 -1484 -38353
rect 1484 -38387 1500 -38353
rect -1500 -38434 1500 -38387
rect -1500 -39481 1500 -39434
rect -1500 -39515 -1484 -39481
rect 1484 -39515 1500 -39481
rect -1500 -39531 1500 -39515
rect -1500 -39589 1500 -39573
rect -1500 -39623 -1484 -39589
rect 1484 -39623 1500 -39589
rect -1500 -39670 1500 -39623
rect -1500 -40717 1500 -40670
rect -1500 -40751 -1484 -40717
rect 1484 -40751 1500 -40717
rect -1500 -40767 1500 -40751
rect -1500 -40825 1500 -40809
rect -1500 -40859 -1484 -40825
rect 1484 -40859 1500 -40825
rect -1500 -40906 1500 -40859
rect -1500 -41953 1500 -41906
rect -1500 -41987 -1484 -41953
rect 1484 -41987 1500 -41953
rect -1500 -42003 1500 -41987
rect -1500 -42061 1500 -42045
rect -1500 -42095 -1484 -42061
rect 1484 -42095 1500 -42061
rect -1500 -42142 1500 -42095
rect -1500 -43189 1500 -43142
rect -1500 -43223 -1484 -43189
rect 1484 -43223 1500 -43189
rect -1500 -43239 1500 -43223
rect -1500 -43297 1500 -43281
rect -1500 -43331 -1484 -43297
rect 1484 -43331 1500 -43297
rect -1500 -43378 1500 -43331
rect -1500 -44425 1500 -44378
rect -1500 -44459 -1484 -44425
rect 1484 -44459 1500 -44425
rect -1500 -44475 1500 -44459
rect -1500 -44533 1500 -44517
rect -1500 -44567 -1484 -44533
rect 1484 -44567 1500 -44533
rect -1500 -44614 1500 -44567
rect -1500 -45661 1500 -45614
rect -1500 -45695 -1484 -45661
rect 1484 -45695 1500 -45661
rect -1500 -45711 1500 -45695
rect -1500 -45769 1500 -45753
rect -1500 -45803 -1484 -45769
rect 1484 -45803 1500 -45769
rect -1500 -45850 1500 -45803
rect -1500 -46897 1500 -46850
rect -1500 -46931 -1484 -46897
rect 1484 -46931 1500 -46897
rect -1500 -46947 1500 -46931
rect -1500 -47005 1500 -46989
rect -1500 -47039 -1484 -47005
rect 1484 -47039 1500 -47005
rect -1500 -47086 1500 -47039
rect -1500 -48133 1500 -48086
rect -1500 -48167 -1484 -48133
rect 1484 -48167 1500 -48133
rect -1500 -48183 1500 -48167
rect -1500 -48241 1500 -48225
rect -1500 -48275 -1484 -48241
rect 1484 -48275 1500 -48241
rect -1500 -48322 1500 -48275
rect -1500 -49369 1500 -49322
rect -1500 -49403 -1484 -49369
rect 1484 -49403 1500 -49369
rect -1500 -49419 1500 -49403
rect -1500 -49477 1500 -49461
rect -1500 -49511 -1484 -49477
rect 1484 -49511 1500 -49477
rect -1500 -49558 1500 -49511
rect -1500 -50605 1500 -50558
rect -1500 -50639 -1484 -50605
rect 1484 -50639 1500 -50605
rect -1500 -50655 1500 -50639
rect -1500 -50713 1500 -50697
rect -1500 -50747 -1484 -50713
rect 1484 -50747 1500 -50713
rect -1500 -50794 1500 -50747
rect -1500 -51841 1500 -51794
rect -1500 -51875 -1484 -51841
rect 1484 -51875 1500 -51841
rect -1500 -51891 1500 -51875
rect -1500 -51949 1500 -51933
rect -1500 -51983 -1484 -51949
rect 1484 -51983 1500 -51949
rect -1500 -52030 1500 -51983
rect -1500 -53077 1500 -53030
rect -1500 -53111 -1484 -53077
rect 1484 -53111 1500 -53077
rect -1500 -53127 1500 -53111
rect -1500 -53185 1500 -53169
rect -1500 -53219 -1484 -53185
rect 1484 -53219 1500 -53185
rect -1500 -53266 1500 -53219
rect -1500 -54313 1500 -54266
rect -1500 -54347 -1484 -54313
rect 1484 -54347 1500 -54313
rect -1500 -54363 1500 -54347
rect -1500 -54421 1500 -54405
rect -1500 -54455 -1484 -54421
rect 1484 -54455 1500 -54421
rect -1500 -54502 1500 -54455
rect -1500 -55549 1500 -55502
rect -1500 -55583 -1484 -55549
rect 1484 -55583 1500 -55549
rect -1500 -55599 1500 -55583
rect -1500 -55657 1500 -55641
rect -1500 -55691 -1484 -55657
rect 1484 -55691 1500 -55657
rect -1500 -55738 1500 -55691
rect -1500 -56785 1500 -56738
rect -1500 -56819 -1484 -56785
rect 1484 -56819 1500 -56785
rect -1500 -56835 1500 -56819
rect -1500 -56893 1500 -56877
rect -1500 -56927 -1484 -56893
rect 1484 -56927 1500 -56893
rect -1500 -56974 1500 -56927
rect -1500 -58021 1500 -57974
rect -1500 -58055 -1484 -58021
rect 1484 -58055 1500 -58021
rect -1500 -58071 1500 -58055
rect -1500 -58129 1500 -58113
rect -1500 -58163 -1484 -58129
rect 1484 -58163 1500 -58129
rect -1500 -58210 1500 -58163
rect -1500 -59257 1500 -59210
rect -1500 -59291 -1484 -59257
rect 1484 -59291 1500 -59257
rect -1500 -59307 1500 -59291
rect -1500 -59365 1500 -59349
rect -1500 -59399 -1484 -59365
rect 1484 -59399 1500 -59365
rect -1500 -59446 1500 -59399
rect -1500 -60493 1500 -60446
rect -1500 -60527 -1484 -60493
rect 1484 -60527 1500 -60493
rect -1500 -60543 1500 -60527
rect -1500 -60601 1500 -60585
rect -1500 -60635 -1484 -60601
rect 1484 -60635 1500 -60601
rect -1500 -60682 1500 -60635
rect -1500 -61729 1500 -61682
rect -1500 -61763 -1484 -61729
rect 1484 -61763 1500 -61729
rect -1500 -61779 1500 -61763
rect -1500 -61837 1500 -61821
rect -1500 -61871 -1484 -61837
rect 1484 -61871 1500 -61837
rect -1500 -61918 1500 -61871
rect -1500 -62965 1500 -62918
rect -1500 -62999 -1484 -62965
rect 1484 -62999 1500 -62965
rect -1500 -63015 1500 -62999
<< polycont >>
rect -1484 62965 1484 62999
rect -1484 61837 1484 61871
rect -1484 61729 1484 61763
rect -1484 60601 1484 60635
rect -1484 60493 1484 60527
rect -1484 59365 1484 59399
rect -1484 59257 1484 59291
rect -1484 58129 1484 58163
rect -1484 58021 1484 58055
rect -1484 56893 1484 56927
rect -1484 56785 1484 56819
rect -1484 55657 1484 55691
rect -1484 55549 1484 55583
rect -1484 54421 1484 54455
rect -1484 54313 1484 54347
rect -1484 53185 1484 53219
rect -1484 53077 1484 53111
rect -1484 51949 1484 51983
rect -1484 51841 1484 51875
rect -1484 50713 1484 50747
rect -1484 50605 1484 50639
rect -1484 49477 1484 49511
rect -1484 49369 1484 49403
rect -1484 48241 1484 48275
rect -1484 48133 1484 48167
rect -1484 47005 1484 47039
rect -1484 46897 1484 46931
rect -1484 45769 1484 45803
rect -1484 45661 1484 45695
rect -1484 44533 1484 44567
rect -1484 44425 1484 44459
rect -1484 43297 1484 43331
rect -1484 43189 1484 43223
rect -1484 42061 1484 42095
rect -1484 41953 1484 41987
rect -1484 40825 1484 40859
rect -1484 40717 1484 40751
rect -1484 39589 1484 39623
rect -1484 39481 1484 39515
rect -1484 38353 1484 38387
rect -1484 38245 1484 38279
rect -1484 37117 1484 37151
rect -1484 37009 1484 37043
rect -1484 35881 1484 35915
rect -1484 35773 1484 35807
rect -1484 34645 1484 34679
rect -1484 34537 1484 34571
rect -1484 33409 1484 33443
rect -1484 33301 1484 33335
rect -1484 32173 1484 32207
rect -1484 32065 1484 32099
rect -1484 30937 1484 30971
rect -1484 30829 1484 30863
rect -1484 29701 1484 29735
rect -1484 29593 1484 29627
rect -1484 28465 1484 28499
rect -1484 28357 1484 28391
rect -1484 27229 1484 27263
rect -1484 27121 1484 27155
rect -1484 25993 1484 26027
rect -1484 25885 1484 25919
rect -1484 24757 1484 24791
rect -1484 24649 1484 24683
rect -1484 23521 1484 23555
rect -1484 23413 1484 23447
rect -1484 22285 1484 22319
rect -1484 22177 1484 22211
rect -1484 21049 1484 21083
rect -1484 20941 1484 20975
rect -1484 19813 1484 19847
rect -1484 19705 1484 19739
rect -1484 18577 1484 18611
rect -1484 18469 1484 18503
rect -1484 17341 1484 17375
rect -1484 17233 1484 17267
rect -1484 16105 1484 16139
rect -1484 15997 1484 16031
rect -1484 14869 1484 14903
rect -1484 14761 1484 14795
rect -1484 13633 1484 13667
rect -1484 13525 1484 13559
rect -1484 12397 1484 12431
rect -1484 12289 1484 12323
rect -1484 11161 1484 11195
rect -1484 11053 1484 11087
rect -1484 9925 1484 9959
rect -1484 9817 1484 9851
rect -1484 8689 1484 8723
rect -1484 8581 1484 8615
rect -1484 7453 1484 7487
rect -1484 7345 1484 7379
rect -1484 6217 1484 6251
rect -1484 6109 1484 6143
rect -1484 4981 1484 5015
rect -1484 4873 1484 4907
rect -1484 3745 1484 3779
rect -1484 3637 1484 3671
rect -1484 2509 1484 2543
rect -1484 2401 1484 2435
rect -1484 1273 1484 1307
rect -1484 1165 1484 1199
rect -1484 37 1484 71
rect -1484 -71 1484 -37
rect -1484 -1199 1484 -1165
rect -1484 -1307 1484 -1273
rect -1484 -2435 1484 -2401
rect -1484 -2543 1484 -2509
rect -1484 -3671 1484 -3637
rect -1484 -3779 1484 -3745
rect -1484 -4907 1484 -4873
rect -1484 -5015 1484 -4981
rect -1484 -6143 1484 -6109
rect -1484 -6251 1484 -6217
rect -1484 -7379 1484 -7345
rect -1484 -7487 1484 -7453
rect -1484 -8615 1484 -8581
rect -1484 -8723 1484 -8689
rect -1484 -9851 1484 -9817
rect -1484 -9959 1484 -9925
rect -1484 -11087 1484 -11053
rect -1484 -11195 1484 -11161
rect -1484 -12323 1484 -12289
rect -1484 -12431 1484 -12397
rect -1484 -13559 1484 -13525
rect -1484 -13667 1484 -13633
rect -1484 -14795 1484 -14761
rect -1484 -14903 1484 -14869
rect -1484 -16031 1484 -15997
rect -1484 -16139 1484 -16105
rect -1484 -17267 1484 -17233
rect -1484 -17375 1484 -17341
rect -1484 -18503 1484 -18469
rect -1484 -18611 1484 -18577
rect -1484 -19739 1484 -19705
rect -1484 -19847 1484 -19813
rect -1484 -20975 1484 -20941
rect -1484 -21083 1484 -21049
rect -1484 -22211 1484 -22177
rect -1484 -22319 1484 -22285
rect -1484 -23447 1484 -23413
rect -1484 -23555 1484 -23521
rect -1484 -24683 1484 -24649
rect -1484 -24791 1484 -24757
rect -1484 -25919 1484 -25885
rect -1484 -26027 1484 -25993
rect -1484 -27155 1484 -27121
rect -1484 -27263 1484 -27229
rect -1484 -28391 1484 -28357
rect -1484 -28499 1484 -28465
rect -1484 -29627 1484 -29593
rect -1484 -29735 1484 -29701
rect -1484 -30863 1484 -30829
rect -1484 -30971 1484 -30937
rect -1484 -32099 1484 -32065
rect -1484 -32207 1484 -32173
rect -1484 -33335 1484 -33301
rect -1484 -33443 1484 -33409
rect -1484 -34571 1484 -34537
rect -1484 -34679 1484 -34645
rect -1484 -35807 1484 -35773
rect -1484 -35915 1484 -35881
rect -1484 -37043 1484 -37009
rect -1484 -37151 1484 -37117
rect -1484 -38279 1484 -38245
rect -1484 -38387 1484 -38353
rect -1484 -39515 1484 -39481
rect -1484 -39623 1484 -39589
rect -1484 -40751 1484 -40717
rect -1484 -40859 1484 -40825
rect -1484 -41987 1484 -41953
rect -1484 -42095 1484 -42061
rect -1484 -43223 1484 -43189
rect -1484 -43331 1484 -43297
rect -1484 -44459 1484 -44425
rect -1484 -44567 1484 -44533
rect -1484 -45695 1484 -45661
rect -1484 -45803 1484 -45769
rect -1484 -46931 1484 -46897
rect -1484 -47039 1484 -47005
rect -1484 -48167 1484 -48133
rect -1484 -48275 1484 -48241
rect -1484 -49403 1484 -49369
rect -1484 -49511 1484 -49477
rect -1484 -50639 1484 -50605
rect -1484 -50747 1484 -50713
rect -1484 -51875 1484 -51841
rect -1484 -51983 1484 -51949
rect -1484 -53111 1484 -53077
rect -1484 -53219 1484 -53185
rect -1484 -54347 1484 -54313
rect -1484 -54455 1484 -54421
rect -1484 -55583 1484 -55549
rect -1484 -55691 1484 -55657
rect -1484 -56819 1484 -56785
rect -1484 -56927 1484 -56893
rect -1484 -58055 1484 -58021
rect -1484 -58163 1484 -58129
rect -1484 -59291 1484 -59257
rect -1484 -59399 1484 -59365
rect -1484 -60527 1484 -60493
rect -1484 -60635 1484 -60601
rect -1484 -61763 1484 -61729
rect -1484 -61871 1484 -61837
rect -1484 -62999 1484 -62965
<< locali >>
rect -1500 62965 -1484 62999
rect 1484 62965 1500 62999
rect -1546 62906 -1512 62922
rect -1546 61914 -1512 61930
rect 1512 62906 1546 62922
rect 1512 61914 1546 61930
rect -1500 61837 -1484 61871
rect 1484 61837 1500 61871
rect -1500 61729 -1484 61763
rect 1484 61729 1500 61763
rect -1546 61670 -1512 61686
rect -1546 60678 -1512 60694
rect 1512 61670 1546 61686
rect 1512 60678 1546 60694
rect -1500 60601 -1484 60635
rect 1484 60601 1500 60635
rect -1500 60493 -1484 60527
rect 1484 60493 1500 60527
rect -1546 60434 -1512 60450
rect -1546 59442 -1512 59458
rect 1512 60434 1546 60450
rect 1512 59442 1546 59458
rect -1500 59365 -1484 59399
rect 1484 59365 1500 59399
rect -1500 59257 -1484 59291
rect 1484 59257 1500 59291
rect -1546 59198 -1512 59214
rect -1546 58206 -1512 58222
rect 1512 59198 1546 59214
rect 1512 58206 1546 58222
rect -1500 58129 -1484 58163
rect 1484 58129 1500 58163
rect -1500 58021 -1484 58055
rect 1484 58021 1500 58055
rect -1546 57962 -1512 57978
rect -1546 56970 -1512 56986
rect 1512 57962 1546 57978
rect 1512 56970 1546 56986
rect -1500 56893 -1484 56927
rect 1484 56893 1500 56927
rect -1500 56785 -1484 56819
rect 1484 56785 1500 56819
rect -1546 56726 -1512 56742
rect -1546 55734 -1512 55750
rect 1512 56726 1546 56742
rect 1512 55734 1546 55750
rect -1500 55657 -1484 55691
rect 1484 55657 1500 55691
rect -1500 55549 -1484 55583
rect 1484 55549 1500 55583
rect -1546 55490 -1512 55506
rect -1546 54498 -1512 54514
rect 1512 55490 1546 55506
rect 1512 54498 1546 54514
rect -1500 54421 -1484 54455
rect 1484 54421 1500 54455
rect -1500 54313 -1484 54347
rect 1484 54313 1500 54347
rect -1546 54254 -1512 54270
rect -1546 53262 -1512 53278
rect 1512 54254 1546 54270
rect 1512 53262 1546 53278
rect -1500 53185 -1484 53219
rect 1484 53185 1500 53219
rect -1500 53077 -1484 53111
rect 1484 53077 1500 53111
rect -1546 53018 -1512 53034
rect -1546 52026 -1512 52042
rect 1512 53018 1546 53034
rect 1512 52026 1546 52042
rect -1500 51949 -1484 51983
rect 1484 51949 1500 51983
rect -1500 51841 -1484 51875
rect 1484 51841 1500 51875
rect -1546 51782 -1512 51798
rect -1546 50790 -1512 50806
rect 1512 51782 1546 51798
rect 1512 50790 1546 50806
rect -1500 50713 -1484 50747
rect 1484 50713 1500 50747
rect -1500 50605 -1484 50639
rect 1484 50605 1500 50639
rect -1546 50546 -1512 50562
rect -1546 49554 -1512 49570
rect 1512 50546 1546 50562
rect 1512 49554 1546 49570
rect -1500 49477 -1484 49511
rect 1484 49477 1500 49511
rect -1500 49369 -1484 49403
rect 1484 49369 1500 49403
rect -1546 49310 -1512 49326
rect -1546 48318 -1512 48334
rect 1512 49310 1546 49326
rect 1512 48318 1546 48334
rect -1500 48241 -1484 48275
rect 1484 48241 1500 48275
rect -1500 48133 -1484 48167
rect 1484 48133 1500 48167
rect -1546 48074 -1512 48090
rect -1546 47082 -1512 47098
rect 1512 48074 1546 48090
rect 1512 47082 1546 47098
rect -1500 47005 -1484 47039
rect 1484 47005 1500 47039
rect -1500 46897 -1484 46931
rect 1484 46897 1500 46931
rect -1546 46838 -1512 46854
rect -1546 45846 -1512 45862
rect 1512 46838 1546 46854
rect 1512 45846 1546 45862
rect -1500 45769 -1484 45803
rect 1484 45769 1500 45803
rect -1500 45661 -1484 45695
rect 1484 45661 1500 45695
rect -1546 45602 -1512 45618
rect -1546 44610 -1512 44626
rect 1512 45602 1546 45618
rect 1512 44610 1546 44626
rect -1500 44533 -1484 44567
rect 1484 44533 1500 44567
rect -1500 44425 -1484 44459
rect 1484 44425 1500 44459
rect -1546 44366 -1512 44382
rect -1546 43374 -1512 43390
rect 1512 44366 1546 44382
rect 1512 43374 1546 43390
rect -1500 43297 -1484 43331
rect 1484 43297 1500 43331
rect -1500 43189 -1484 43223
rect 1484 43189 1500 43223
rect -1546 43130 -1512 43146
rect -1546 42138 -1512 42154
rect 1512 43130 1546 43146
rect 1512 42138 1546 42154
rect -1500 42061 -1484 42095
rect 1484 42061 1500 42095
rect -1500 41953 -1484 41987
rect 1484 41953 1500 41987
rect -1546 41894 -1512 41910
rect -1546 40902 -1512 40918
rect 1512 41894 1546 41910
rect 1512 40902 1546 40918
rect -1500 40825 -1484 40859
rect 1484 40825 1500 40859
rect -1500 40717 -1484 40751
rect 1484 40717 1500 40751
rect -1546 40658 -1512 40674
rect -1546 39666 -1512 39682
rect 1512 40658 1546 40674
rect 1512 39666 1546 39682
rect -1500 39589 -1484 39623
rect 1484 39589 1500 39623
rect -1500 39481 -1484 39515
rect 1484 39481 1500 39515
rect -1546 39422 -1512 39438
rect -1546 38430 -1512 38446
rect 1512 39422 1546 39438
rect 1512 38430 1546 38446
rect -1500 38353 -1484 38387
rect 1484 38353 1500 38387
rect -1500 38245 -1484 38279
rect 1484 38245 1500 38279
rect -1546 38186 -1512 38202
rect -1546 37194 -1512 37210
rect 1512 38186 1546 38202
rect 1512 37194 1546 37210
rect -1500 37117 -1484 37151
rect 1484 37117 1500 37151
rect -1500 37009 -1484 37043
rect 1484 37009 1500 37043
rect -1546 36950 -1512 36966
rect -1546 35958 -1512 35974
rect 1512 36950 1546 36966
rect 1512 35958 1546 35974
rect -1500 35881 -1484 35915
rect 1484 35881 1500 35915
rect -1500 35773 -1484 35807
rect 1484 35773 1500 35807
rect -1546 35714 -1512 35730
rect -1546 34722 -1512 34738
rect 1512 35714 1546 35730
rect 1512 34722 1546 34738
rect -1500 34645 -1484 34679
rect 1484 34645 1500 34679
rect -1500 34537 -1484 34571
rect 1484 34537 1500 34571
rect -1546 34478 -1512 34494
rect -1546 33486 -1512 33502
rect 1512 34478 1546 34494
rect 1512 33486 1546 33502
rect -1500 33409 -1484 33443
rect 1484 33409 1500 33443
rect -1500 33301 -1484 33335
rect 1484 33301 1500 33335
rect -1546 33242 -1512 33258
rect -1546 32250 -1512 32266
rect 1512 33242 1546 33258
rect 1512 32250 1546 32266
rect -1500 32173 -1484 32207
rect 1484 32173 1500 32207
rect -1500 32065 -1484 32099
rect 1484 32065 1500 32099
rect -1546 32006 -1512 32022
rect -1546 31014 -1512 31030
rect 1512 32006 1546 32022
rect 1512 31014 1546 31030
rect -1500 30937 -1484 30971
rect 1484 30937 1500 30971
rect -1500 30829 -1484 30863
rect 1484 30829 1500 30863
rect -1546 30770 -1512 30786
rect -1546 29778 -1512 29794
rect 1512 30770 1546 30786
rect 1512 29778 1546 29794
rect -1500 29701 -1484 29735
rect 1484 29701 1500 29735
rect -1500 29593 -1484 29627
rect 1484 29593 1500 29627
rect -1546 29534 -1512 29550
rect -1546 28542 -1512 28558
rect 1512 29534 1546 29550
rect 1512 28542 1546 28558
rect -1500 28465 -1484 28499
rect 1484 28465 1500 28499
rect -1500 28357 -1484 28391
rect 1484 28357 1500 28391
rect -1546 28298 -1512 28314
rect -1546 27306 -1512 27322
rect 1512 28298 1546 28314
rect 1512 27306 1546 27322
rect -1500 27229 -1484 27263
rect 1484 27229 1500 27263
rect -1500 27121 -1484 27155
rect 1484 27121 1500 27155
rect -1546 27062 -1512 27078
rect -1546 26070 -1512 26086
rect 1512 27062 1546 27078
rect 1512 26070 1546 26086
rect -1500 25993 -1484 26027
rect 1484 25993 1500 26027
rect -1500 25885 -1484 25919
rect 1484 25885 1500 25919
rect -1546 25826 -1512 25842
rect -1546 24834 -1512 24850
rect 1512 25826 1546 25842
rect 1512 24834 1546 24850
rect -1500 24757 -1484 24791
rect 1484 24757 1500 24791
rect -1500 24649 -1484 24683
rect 1484 24649 1500 24683
rect -1546 24590 -1512 24606
rect -1546 23598 -1512 23614
rect 1512 24590 1546 24606
rect 1512 23598 1546 23614
rect -1500 23521 -1484 23555
rect 1484 23521 1500 23555
rect -1500 23413 -1484 23447
rect 1484 23413 1500 23447
rect -1546 23354 -1512 23370
rect -1546 22362 -1512 22378
rect 1512 23354 1546 23370
rect 1512 22362 1546 22378
rect -1500 22285 -1484 22319
rect 1484 22285 1500 22319
rect -1500 22177 -1484 22211
rect 1484 22177 1500 22211
rect -1546 22118 -1512 22134
rect -1546 21126 -1512 21142
rect 1512 22118 1546 22134
rect 1512 21126 1546 21142
rect -1500 21049 -1484 21083
rect 1484 21049 1500 21083
rect -1500 20941 -1484 20975
rect 1484 20941 1500 20975
rect -1546 20882 -1512 20898
rect -1546 19890 -1512 19906
rect 1512 20882 1546 20898
rect 1512 19890 1546 19906
rect -1500 19813 -1484 19847
rect 1484 19813 1500 19847
rect -1500 19705 -1484 19739
rect 1484 19705 1500 19739
rect -1546 19646 -1512 19662
rect -1546 18654 -1512 18670
rect 1512 19646 1546 19662
rect 1512 18654 1546 18670
rect -1500 18577 -1484 18611
rect 1484 18577 1500 18611
rect -1500 18469 -1484 18503
rect 1484 18469 1500 18503
rect -1546 18410 -1512 18426
rect -1546 17418 -1512 17434
rect 1512 18410 1546 18426
rect 1512 17418 1546 17434
rect -1500 17341 -1484 17375
rect 1484 17341 1500 17375
rect -1500 17233 -1484 17267
rect 1484 17233 1500 17267
rect -1546 17174 -1512 17190
rect -1546 16182 -1512 16198
rect 1512 17174 1546 17190
rect 1512 16182 1546 16198
rect -1500 16105 -1484 16139
rect 1484 16105 1500 16139
rect -1500 15997 -1484 16031
rect 1484 15997 1500 16031
rect -1546 15938 -1512 15954
rect -1546 14946 -1512 14962
rect 1512 15938 1546 15954
rect 1512 14946 1546 14962
rect -1500 14869 -1484 14903
rect 1484 14869 1500 14903
rect -1500 14761 -1484 14795
rect 1484 14761 1500 14795
rect -1546 14702 -1512 14718
rect -1546 13710 -1512 13726
rect 1512 14702 1546 14718
rect 1512 13710 1546 13726
rect -1500 13633 -1484 13667
rect 1484 13633 1500 13667
rect -1500 13525 -1484 13559
rect 1484 13525 1500 13559
rect -1546 13466 -1512 13482
rect -1546 12474 -1512 12490
rect 1512 13466 1546 13482
rect 1512 12474 1546 12490
rect -1500 12397 -1484 12431
rect 1484 12397 1500 12431
rect -1500 12289 -1484 12323
rect 1484 12289 1500 12323
rect -1546 12230 -1512 12246
rect -1546 11238 -1512 11254
rect 1512 12230 1546 12246
rect 1512 11238 1546 11254
rect -1500 11161 -1484 11195
rect 1484 11161 1500 11195
rect -1500 11053 -1484 11087
rect 1484 11053 1500 11087
rect -1546 10994 -1512 11010
rect -1546 10002 -1512 10018
rect 1512 10994 1546 11010
rect 1512 10002 1546 10018
rect -1500 9925 -1484 9959
rect 1484 9925 1500 9959
rect -1500 9817 -1484 9851
rect 1484 9817 1500 9851
rect -1546 9758 -1512 9774
rect -1546 8766 -1512 8782
rect 1512 9758 1546 9774
rect 1512 8766 1546 8782
rect -1500 8689 -1484 8723
rect 1484 8689 1500 8723
rect -1500 8581 -1484 8615
rect 1484 8581 1500 8615
rect -1546 8522 -1512 8538
rect -1546 7530 -1512 7546
rect 1512 8522 1546 8538
rect 1512 7530 1546 7546
rect -1500 7453 -1484 7487
rect 1484 7453 1500 7487
rect -1500 7345 -1484 7379
rect 1484 7345 1500 7379
rect -1546 7286 -1512 7302
rect -1546 6294 -1512 6310
rect 1512 7286 1546 7302
rect 1512 6294 1546 6310
rect -1500 6217 -1484 6251
rect 1484 6217 1500 6251
rect -1500 6109 -1484 6143
rect 1484 6109 1500 6143
rect -1546 6050 -1512 6066
rect -1546 5058 -1512 5074
rect 1512 6050 1546 6066
rect 1512 5058 1546 5074
rect -1500 4981 -1484 5015
rect 1484 4981 1500 5015
rect -1500 4873 -1484 4907
rect 1484 4873 1500 4907
rect -1546 4814 -1512 4830
rect -1546 3822 -1512 3838
rect 1512 4814 1546 4830
rect 1512 3822 1546 3838
rect -1500 3745 -1484 3779
rect 1484 3745 1500 3779
rect -1500 3637 -1484 3671
rect 1484 3637 1500 3671
rect -1546 3578 -1512 3594
rect -1546 2586 -1512 2602
rect 1512 3578 1546 3594
rect 1512 2586 1546 2602
rect -1500 2509 -1484 2543
rect 1484 2509 1500 2543
rect -1500 2401 -1484 2435
rect 1484 2401 1500 2435
rect -1546 2342 -1512 2358
rect -1546 1350 -1512 1366
rect 1512 2342 1546 2358
rect 1512 1350 1546 1366
rect -1500 1273 -1484 1307
rect 1484 1273 1500 1307
rect -1500 1165 -1484 1199
rect 1484 1165 1500 1199
rect -1546 1106 -1512 1122
rect -1546 114 -1512 130
rect 1512 1106 1546 1122
rect 1512 114 1546 130
rect -1500 37 -1484 71
rect 1484 37 1500 71
rect -1500 -71 -1484 -37
rect 1484 -71 1500 -37
rect -1546 -130 -1512 -114
rect -1546 -1122 -1512 -1106
rect 1512 -130 1546 -114
rect 1512 -1122 1546 -1106
rect -1500 -1199 -1484 -1165
rect 1484 -1199 1500 -1165
rect -1500 -1307 -1484 -1273
rect 1484 -1307 1500 -1273
rect -1546 -1366 -1512 -1350
rect -1546 -2358 -1512 -2342
rect 1512 -1366 1546 -1350
rect 1512 -2358 1546 -2342
rect -1500 -2435 -1484 -2401
rect 1484 -2435 1500 -2401
rect -1500 -2543 -1484 -2509
rect 1484 -2543 1500 -2509
rect -1546 -2602 -1512 -2586
rect -1546 -3594 -1512 -3578
rect 1512 -2602 1546 -2586
rect 1512 -3594 1546 -3578
rect -1500 -3671 -1484 -3637
rect 1484 -3671 1500 -3637
rect -1500 -3779 -1484 -3745
rect 1484 -3779 1500 -3745
rect -1546 -3838 -1512 -3822
rect -1546 -4830 -1512 -4814
rect 1512 -3838 1546 -3822
rect 1512 -4830 1546 -4814
rect -1500 -4907 -1484 -4873
rect 1484 -4907 1500 -4873
rect -1500 -5015 -1484 -4981
rect 1484 -5015 1500 -4981
rect -1546 -5074 -1512 -5058
rect -1546 -6066 -1512 -6050
rect 1512 -5074 1546 -5058
rect 1512 -6066 1546 -6050
rect -1500 -6143 -1484 -6109
rect 1484 -6143 1500 -6109
rect -1500 -6251 -1484 -6217
rect 1484 -6251 1500 -6217
rect -1546 -6310 -1512 -6294
rect -1546 -7302 -1512 -7286
rect 1512 -6310 1546 -6294
rect 1512 -7302 1546 -7286
rect -1500 -7379 -1484 -7345
rect 1484 -7379 1500 -7345
rect -1500 -7487 -1484 -7453
rect 1484 -7487 1500 -7453
rect -1546 -7546 -1512 -7530
rect -1546 -8538 -1512 -8522
rect 1512 -7546 1546 -7530
rect 1512 -8538 1546 -8522
rect -1500 -8615 -1484 -8581
rect 1484 -8615 1500 -8581
rect -1500 -8723 -1484 -8689
rect 1484 -8723 1500 -8689
rect -1546 -8782 -1512 -8766
rect -1546 -9774 -1512 -9758
rect 1512 -8782 1546 -8766
rect 1512 -9774 1546 -9758
rect -1500 -9851 -1484 -9817
rect 1484 -9851 1500 -9817
rect -1500 -9959 -1484 -9925
rect 1484 -9959 1500 -9925
rect -1546 -10018 -1512 -10002
rect -1546 -11010 -1512 -10994
rect 1512 -10018 1546 -10002
rect 1512 -11010 1546 -10994
rect -1500 -11087 -1484 -11053
rect 1484 -11087 1500 -11053
rect -1500 -11195 -1484 -11161
rect 1484 -11195 1500 -11161
rect -1546 -11254 -1512 -11238
rect -1546 -12246 -1512 -12230
rect 1512 -11254 1546 -11238
rect 1512 -12246 1546 -12230
rect -1500 -12323 -1484 -12289
rect 1484 -12323 1500 -12289
rect -1500 -12431 -1484 -12397
rect 1484 -12431 1500 -12397
rect -1546 -12490 -1512 -12474
rect -1546 -13482 -1512 -13466
rect 1512 -12490 1546 -12474
rect 1512 -13482 1546 -13466
rect -1500 -13559 -1484 -13525
rect 1484 -13559 1500 -13525
rect -1500 -13667 -1484 -13633
rect 1484 -13667 1500 -13633
rect -1546 -13726 -1512 -13710
rect -1546 -14718 -1512 -14702
rect 1512 -13726 1546 -13710
rect 1512 -14718 1546 -14702
rect -1500 -14795 -1484 -14761
rect 1484 -14795 1500 -14761
rect -1500 -14903 -1484 -14869
rect 1484 -14903 1500 -14869
rect -1546 -14962 -1512 -14946
rect -1546 -15954 -1512 -15938
rect 1512 -14962 1546 -14946
rect 1512 -15954 1546 -15938
rect -1500 -16031 -1484 -15997
rect 1484 -16031 1500 -15997
rect -1500 -16139 -1484 -16105
rect 1484 -16139 1500 -16105
rect -1546 -16198 -1512 -16182
rect -1546 -17190 -1512 -17174
rect 1512 -16198 1546 -16182
rect 1512 -17190 1546 -17174
rect -1500 -17267 -1484 -17233
rect 1484 -17267 1500 -17233
rect -1500 -17375 -1484 -17341
rect 1484 -17375 1500 -17341
rect -1546 -17434 -1512 -17418
rect -1546 -18426 -1512 -18410
rect 1512 -17434 1546 -17418
rect 1512 -18426 1546 -18410
rect -1500 -18503 -1484 -18469
rect 1484 -18503 1500 -18469
rect -1500 -18611 -1484 -18577
rect 1484 -18611 1500 -18577
rect -1546 -18670 -1512 -18654
rect -1546 -19662 -1512 -19646
rect 1512 -18670 1546 -18654
rect 1512 -19662 1546 -19646
rect -1500 -19739 -1484 -19705
rect 1484 -19739 1500 -19705
rect -1500 -19847 -1484 -19813
rect 1484 -19847 1500 -19813
rect -1546 -19906 -1512 -19890
rect -1546 -20898 -1512 -20882
rect 1512 -19906 1546 -19890
rect 1512 -20898 1546 -20882
rect -1500 -20975 -1484 -20941
rect 1484 -20975 1500 -20941
rect -1500 -21083 -1484 -21049
rect 1484 -21083 1500 -21049
rect -1546 -21142 -1512 -21126
rect -1546 -22134 -1512 -22118
rect 1512 -21142 1546 -21126
rect 1512 -22134 1546 -22118
rect -1500 -22211 -1484 -22177
rect 1484 -22211 1500 -22177
rect -1500 -22319 -1484 -22285
rect 1484 -22319 1500 -22285
rect -1546 -22378 -1512 -22362
rect -1546 -23370 -1512 -23354
rect 1512 -22378 1546 -22362
rect 1512 -23370 1546 -23354
rect -1500 -23447 -1484 -23413
rect 1484 -23447 1500 -23413
rect -1500 -23555 -1484 -23521
rect 1484 -23555 1500 -23521
rect -1546 -23614 -1512 -23598
rect -1546 -24606 -1512 -24590
rect 1512 -23614 1546 -23598
rect 1512 -24606 1546 -24590
rect -1500 -24683 -1484 -24649
rect 1484 -24683 1500 -24649
rect -1500 -24791 -1484 -24757
rect 1484 -24791 1500 -24757
rect -1546 -24850 -1512 -24834
rect -1546 -25842 -1512 -25826
rect 1512 -24850 1546 -24834
rect 1512 -25842 1546 -25826
rect -1500 -25919 -1484 -25885
rect 1484 -25919 1500 -25885
rect -1500 -26027 -1484 -25993
rect 1484 -26027 1500 -25993
rect -1546 -26086 -1512 -26070
rect -1546 -27078 -1512 -27062
rect 1512 -26086 1546 -26070
rect 1512 -27078 1546 -27062
rect -1500 -27155 -1484 -27121
rect 1484 -27155 1500 -27121
rect -1500 -27263 -1484 -27229
rect 1484 -27263 1500 -27229
rect -1546 -27322 -1512 -27306
rect -1546 -28314 -1512 -28298
rect 1512 -27322 1546 -27306
rect 1512 -28314 1546 -28298
rect -1500 -28391 -1484 -28357
rect 1484 -28391 1500 -28357
rect -1500 -28499 -1484 -28465
rect 1484 -28499 1500 -28465
rect -1546 -28558 -1512 -28542
rect -1546 -29550 -1512 -29534
rect 1512 -28558 1546 -28542
rect 1512 -29550 1546 -29534
rect -1500 -29627 -1484 -29593
rect 1484 -29627 1500 -29593
rect -1500 -29735 -1484 -29701
rect 1484 -29735 1500 -29701
rect -1546 -29794 -1512 -29778
rect -1546 -30786 -1512 -30770
rect 1512 -29794 1546 -29778
rect 1512 -30786 1546 -30770
rect -1500 -30863 -1484 -30829
rect 1484 -30863 1500 -30829
rect -1500 -30971 -1484 -30937
rect 1484 -30971 1500 -30937
rect -1546 -31030 -1512 -31014
rect -1546 -32022 -1512 -32006
rect 1512 -31030 1546 -31014
rect 1512 -32022 1546 -32006
rect -1500 -32099 -1484 -32065
rect 1484 -32099 1500 -32065
rect -1500 -32207 -1484 -32173
rect 1484 -32207 1500 -32173
rect -1546 -32266 -1512 -32250
rect -1546 -33258 -1512 -33242
rect 1512 -32266 1546 -32250
rect 1512 -33258 1546 -33242
rect -1500 -33335 -1484 -33301
rect 1484 -33335 1500 -33301
rect -1500 -33443 -1484 -33409
rect 1484 -33443 1500 -33409
rect -1546 -33502 -1512 -33486
rect -1546 -34494 -1512 -34478
rect 1512 -33502 1546 -33486
rect 1512 -34494 1546 -34478
rect -1500 -34571 -1484 -34537
rect 1484 -34571 1500 -34537
rect -1500 -34679 -1484 -34645
rect 1484 -34679 1500 -34645
rect -1546 -34738 -1512 -34722
rect -1546 -35730 -1512 -35714
rect 1512 -34738 1546 -34722
rect 1512 -35730 1546 -35714
rect -1500 -35807 -1484 -35773
rect 1484 -35807 1500 -35773
rect -1500 -35915 -1484 -35881
rect 1484 -35915 1500 -35881
rect -1546 -35974 -1512 -35958
rect -1546 -36966 -1512 -36950
rect 1512 -35974 1546 -35958
rect 1512 -36966 1546 -36950
rect -1500 -37043 -1484 -37009
rect 1484 -37043 1500 -37009
rect -1500 -37151 -1484 -37117
rect 1484 -37151 1500 -37117
rect -1546 -37210 -1512 -37194
rect -1546 -38202 -1512 -38186
rect 1512 -37210 1546 -37194
rect 1512 -38202 1546 -38186
rect -1500 -38279 -1484 -38245
rect 1484 -38279 1500 -38245
rect -1500 -38387 -1484 -38353
rect 1484 -38387 1500 -38353
rect -1546 -38446 -1512 -38430
rect -1546 -39438 -1512 -39422
rect 1512 -38446 1546 -38430
rect 1512 -39438 1546 -39422
rect -1500 -39515 -1484 -39481
rect 1484 -39515 1500 -39481
rect -1500 -39623 -1484 -39589
rect 1484 -39623 1500 -39589
rect -1546 -39682 -1512 -39666
rect -1546 -40674 -1512 -40658
rect 1512 -39682 1546 -39666
rect 1512 -40674 1546 -40658
rect -1500 -40751 -1484 -40717
rect 1484 -40751 1500 -40717
rect -1500 -40859 -1484 -40825
rect 1484 -40859 1500 -40825
rect -1546 -40918 -1512 -40902
rect -1546 -41910 -1512 -41894
rect 1512 -40918 1546 -40902
rect 1512 -41910 1546 -41894
rect -1500 -41987 -1484 -41953
rect 1484 -41987 1500 -41953
rect -1500 -42095 -1484 -42061
rect 1484 -42095 1500 -42061
rect -1546 -42154 -1512 -42138
rect -1546 -43146 -1512 -43130
rect 1512 -42154 1546 -42138
rect 1512 -43146 1546 -43130
rect -1500 -43223 -1484 -43189
rect 1484 -43223 1500 -43189
rect -1500 -43331 -1484 -43297
rect 1484 -43331 1500 -43297
rect -1546 -43390 -1512 -43374
rect -1546 -44382 -1512 -44366
rect 1512 -43390 1546 -43374
rect 1512 -44382 1546 -44366
rect -1500 -44459 -1484 -44425
rect 1484 -44459 1500 -44425
rect -1500 -44567 -1484 -44533
rect 1484 -44567 1500 -44533
rect -1546 -44626 -1512 -44610
rect -1546 -45618 -1512 -45602
rect 1512 -44626 1546 -44610
rect 1512 -45618 1546 -45602
rect -1500 -45695 -1484 -45661
rect 1484 -45695 1500 -45661
rect -1500 -45803 -1484 -45769
rect 1484 -45803 1500 -45769
rect -1546 -45862 -1512 -45846
rect -1546 -46854 -1512 -46838
rect 1512 -45862 1546 -45846
rect 1512 -46854 1546 -46838
rect -1500 -46931 -1484 -46897
rect 1484 -46931 1500 -46897
rect -1500 -47039 -1484 -47005
rect 1484 -47039 1500 -47005
rect -1546 -47098 -1512 -47082
rect -1546 -48090 -1512 -48074
rect 1512 -47098 1546 -47082
rect 1512 -48090 1546 -48074
rect -1500 -48167 -1484 -48133
rect 1484 -48167 1500 -48133
rect -1500 -48275 -1484 -48241
rect 1484 -48275 1500 -48241
rect -1546 -48334 -1512 -48318
rect -1546 -49326 -1512 -49310
rect 1512 -48334 1546 -48318
rect 1512 -49326 1546 -49310
rect -1500 -49403 -1484 -49369
rect 1484 -49403 1500 -49369
rect -1500 -49511 -1484 -49477
rect 1484 -49511 1500 -49477
rect -1546 -49570 -1512 -49554
rect -1546 -50562 -1512 -50546
rect 1512 -49570 1546 -49554
rect 1512 -50562 1546 -50546
rect -1500 -50639 -1484 -50605
rect 1484 -50639 1500 -50605
rect -1500 -50747 -1484 -50713
rect 1484 -50747 1500 -50713
rect -1546 -50806 -1512 -50790
rect -1546 -51798 -1512 -51782
rect 1512 -50806 1546 -50790
rect 1512 -51798 1546 -51782
rect -1500 -51875 -1484 -51841
rect 1484 -51875 1500 -51841
rect -1500 -51983 -1484 -51949
rect 1484 -51983 1500 -51949
rect -1546 -52042 -1512 -52026
rect -1546 -53034 -1512 -53018
rect 1512 -52042 1546 -52026
rect 1512 -53034 1546 -53018
rect -1500 -53111 -1484 -53077
rect 1484 -53111 1500 -53077
rect -1500 -53219 -1484 -53185
rect 1484 -53219 1500 -53185
rect -1546 -53278 -1512 -53262
rect -1546 -54270 -1512 -54254
rect 1512 -53278 1546 -53262
rect 1512 -54270 1546 -54254
rect -1500 -54347 -1484 -54313
rect 1484 -54347 1500 -54313
rect -1500 -54455 -1484 -54421
rect 1484 -54455 1500 -54421
rect -1546 -54514 -1512 -54498
rect -1546 -55506 -1512 -55490
rect 1512 -54514 1546 -54498
rect 1512 -55506 1546 -55490
rect -1500 -55583 -1484 -55549
rect 1484 -55583 1500 -55549
rect -1500 -55691 -1484 -55657
rect 1484 -55691 1500 -55657
rect -1546 -55750 -1512 -55734
rect -1546 -56742 -1512 -56726
rect 1512 -55750 1546 -55734
rect 1512 -56742 1546 -56726
rect -1500 -56819 -1484 -56785
rect 1484 -56819 1500 -56785
rect -1500 -56927 -1484 -56893
rect 1484 -56927 1500 -56893
rect -1546 -56986 -1512 -56970
rect -1546 -57978 -1512 -57962
rect 1512 -56986 1546 -56970
rect 1512 -57978 1546 -57962
rect -1500 -58055 -1484 -58021
rect 1484 -58055 1500 -58021
rect -1500 -58163 -1484 -58129
rect 1484 -58163 1500 -58129
rect -1546 -58222 -1512 -58206
rect -1546 -59214 -1512 -59198
rect 1512 -58222 1546 -58206
rect 1512 -59214 1546 -59198
rect -1500 -59291 -1484 -59257
rect 1484 -59291 1500 -59257
rect -1500 -59399 -1484 -59365
rect 1484 -59399 1500 -59365
rect -1546 -59458 -1512 -59442
rect -1546 -60450 -1512 -60434
rect 1512 -59458 1546 -59442
rect 1512 -60450 1546 -60434
rect -1500 -60527 -1484 -60493
rect 1484 -60527 1500 -60493
rect -1500 -60635 -1484 -60601
rect 1484 -60635 1500 -60601
rect -1546 -60694 -1512 -60678
rect -1546 -61686 -1512 -61670
rect 1512 -60694 1546 -60678
rect 1512 -61686 1546 -61670
rect -1500 -61763 -1484 -61729
rect 1484 -61763 1500 -61729
rect -1500 -61871 -1484 -61837
rect 1484 -61871 1500 -61837
rect -1546 -61930 -1512 -61914
rect -1546 -62922 -1512 -62906
rect 1512 -61930 1546 -61914
rect 1512 -62922 1546 -62906
rect -1500 -62999 -1484 -62965
rect 1484 -62999 1500 -62965
<< viali >>
rect -1484 62965 1484 62999
rect -1546 61930 -1512 62906
rect 1512 61930 1546 62906
rect -1484 61837 1484 61871
rect -1484 61729 1484 61763
rect -1546 60694 -1512 61670
rect 1512 60694 1546 61670
rect -1484 60601 1484 60635
rect -1484 60493 1484 60527
rect -1546 59458 -1512 60434
rect 1512 59458 1546 60434
rect -1484 59365 1484 59399
rect -1484 59257 1484 59291
rect -1546 58222 -1512 59198
rect 1512 58222 1546 59198
rect -1484 58129 1484 58163
rect -1484 58021 1484 58055
rect -1546 56986 -1512 57962
rect 1512 56986 1546 57962
rect -1484 56893 1484 56927
rect -1484 56785 1484 56819
rect -1546 55750 -1512 56726
rect 1512 55750 1546 56726
rect -1484 55657 1484 55691
rect -1484 55549 1484 55583
rect -1546 54514 -1512 55490
rect 1512 54514 1546 55490
rect -1484 54421 1484 54455
rect -1484 54313 1484 54347
rect -1546 53278 -1512 54254
rect 1512 53278 1546 54254
rect -1484 53185 1484 53219
rect -1484 53077 1484 53111
rect -1546 52042 -1512 53018
rect 1512 52042 1546 53018
rect -1484 51949 1484 51983
rect -1484 51841 1484 51875
rect -1546 50806 -1512 51782
rect 1512 50806 1546 51782
rect -1484 50713 1484 50747
rect -1484 50605 1484 50639
rect -1546 49570 -1512 50546
rect 1512 49570 1546 50546
rect -1484 49477 1484 49511
rect -1484 49369 1484 49403
rect -1546 48334 -1512 49310
rect 1512 48334 1546 49310
rect -1484 48241 1484 48275
rect -1484 48133 1484 48167
rect -1546 47098 -1512 48074
rect 1512 47098 1546 48074
rect -1484 47005 1484 47039
rect -1484 46897 1484 46931
rect -1546 45862 -1512 46838
rect 1512 45862 1546 46838
rect -1484 45769 1484 45803
rect -1484 45661 1484 45695
rect -1546 44626 -1512 45602
rect 1512 44626 1546 45602
rect -1484 44533 1484 44567
rect -1484 44425 1484 44459
rect -1546 43390 -1512 44366
rect 1512 43390 1546 44366
rect -1484 43297 1484 43331
rect -1484 43189 1484 43223
rect -1546 42154 -1512 43130
rect 1512 42154 1546 43130
rect -1484 42061 1484 42095
rect -1484 41953 1484 41987
rect -1546 40918 -1512 41894
rect 1512 40918 1546 41894
rect -1484 40825 1484 40859
rect -1484 40717 1484 40751
rect -1546 39682 -1512 40658
rect 1512 39682 1546 40658
rect -1484 39589 1484 39623
rect -1484 39481 1484 39515
rect -1546 38446 -1512 39422
rect 1512 38446 1546 39422
rect -1484 38353 1484 38387
rect -1484 38245 1484 38279
rect -1546 37210 -1512 38186
rect 1512 37210 1546 38186
rect -1484 37117 1484 37151
rect -1484 37009 1484 37043
rect -1546 35974 -1512 36950
rect 1512 35974 1546 36950
rect -1484 35881 1484 35915
rect -1484 35773 1484 35807
rect -1546 34738 -1512 35714
rect 1512 34738 1546 35714
rect -1484 34645 1484 34679
rect -1484 34537 1484 34571
rect -1546 33502 -1512 34478
rect 1512 33502 1546 34478
rect -1484 33409 1484 33443
rect -1484 33301 1484 33335
rect -1546 32266 -1512 33242
rect 1512 32266 1546 33242
rect -1484 32173 1484 32207
rect -1484 32065 1484 32099
rect -1546 31030 -1512 32006
rect 1512 31030 1546 32006
rect -1484 30937 1484 30971
rect -1484 30829 1484 30863
rect -1546 29794 -1512 30770
rect 1512 29794 1546 30770
rect -1484 29701 1484 29735
rect -1484 29593 1484 29627
rect -1546 28558 -1512 29534
rect 1512 28558 1546 29534
rect -1484 28465 1484 28499
rect -1484 28357 1484 28391
rect -1546 27322 -1512 28298
rect 1512 27322 1546 28298
rect -1484 27229 1484 27263
rect -1484 27121 1484 27155
rect -1546 26086 -1512 27062
rect 1512 26086 1546 27062
rect -1484 25993 1484 26027
rect -1484 25885 1484 25919
rect -1546 24850 -1512 25826
rect 1512 24850 1546 25826
rect -1484 24757 1484 24791
rect -1484 24649 1484 24683
rect -1546 23614 -1512 24590
rect 1512 23614 1546 24590
rect -1484 23521 1484 23555
rect -1484 23413 1484 23447
rect -1546 22378 -1512 23354
rect 1512 22378 1546 23354
rect -1484 22285 1484 22319
rect -1484 22177 1484 22211
rect -1546 21142 -1512 22118
rect 1512 21142 1546 22118
rect -1484 21049 1484 21083
rect -1484 20941 1484 20975
rect -1546 19906 -1512 20882
rect 1512 19906 1546 20882
rect -1484 19813 1484 19847
rect -1484 19705 1484 19739
rect -1546 18670 -1512 19646
rect 1512 18670 1546 19646
rect -1484 18577 1484 18611
rect -1484 18469 1484 18503
rect -1546 17434 -1512 18410
rect 1512 17434 1546 18410
rect -1484 17341 1484 17375
rect -1484 17233 1484 17267
rect -1546 16198 -1512 17174
rect 1512 16198 1546 17174
rect -1484 16105 1484 16139
rect -1484 15997 1484 16031
rect -1546 14962 -1512 15938
rect 1512 14962 1546 15938
rect -1484 14869 1484 14903
rect -1484 14761 1484 14795
rect -1546 13726 -1512 14702
rect 1512 13726 1546 14702
rect -1484 13633 1484 13667
rect -1484 13525 1484 13559
rect -1546 12490 -1512 13466
rect 1512 12490 1546 13466
rect -1484 12397 1484 12431
rect -1484 12289 1484 12323
rect -1546 11254 -1512 12230
rect 1512 11254 1546 12230
rect -1484 11161 1484 11195
rect -1484 11053 1484 11087
rect -1546 10018 -1512 10994
rect 1512 10018 1546 10994
rect -1484 9925 1484 9959
rect -1484 9817 1484 9851
rect -1546 8782 -1512 9758
rect 1512 8782 1546 9758
rect -1484 8689 1484 8723
rect -1484 8581 1484 8615
rect -1546 7546 -1512 8522
rect 1512 7546 1546 8522
rect -1484 7453 1484 7487
rect -1484 7345 1484 7379
rect -1546 6310 -1512 7286
rect 1512 6310 1546 7286
rect -1484 6217 1484 6251
rect -1484 6109 1484 6143
rect -1546 5074 -1512 6050
rect 1512 5074 1546 6050
rect -1484 4981 1484 5015
rect -1484 4873 1484 4907
rect -1546 3838 -1512 4814
rect 1512 3838 1546 4814
rect -1484 3745 1484 3779
rect -1484 3637 1484 3671
rect -1546 2602 -1512 3578
rect 1512 2602 1546 3578
rect -1484 2509 1484 2543
rect -1484 2401 1484 2435
rect -1546 1366 -1512 2342
rect 1512 1366 1546 2342
rect -1484 1273 1484 1307
rect -1484 1165 1484 1199
rect -1546 130 -1512 1106
rect 1512 130 1546 1106
rect -1484 37 1484 71
rect -1484 -71 1484 -37
rect -1546 -1106 -1512 -130
rect 1512 -1106 1546 -130
rect -1484 -1199 1484 -1165
rect -1484 -1307 1484 -1273
rect -1546 -2342 -1512 -1366
rect 1512 -2342 1546 -1366
rect -1484 -2435 1484 -2401
rect -1484 -2543 1484 -2509
rect -1546 -3578 -1512 -2602
rect 1512 -3578 1546 -2602
rect -1484 -3671 1484 -3637
rect -1484 -3779 1484 -3745
rect -1546 -4814 -1512 -3838
rect 1512 -4814 1546 -3838
rect -1484 -4907 1484 -4873
rect -1484 -5015 1484 -4981
rect -1546 -6050 -1512 -5074
rect 1512 -6050 1546 -5074
rect -1484 -6143 1484 -6109
rect -1484 -6251 1484 -6217
rect -1546 -7286 -1512 -6310
rect 1512 -7286 1546 -6310
rect -1484 -7379 1484 -7345
rect -1484 -7487 1484 -7453
rect -1546 -8522 -1512 -7546
rect 1512 -8522 1546 -7546
rect -1484 -8615 1484 -8581
rect -1484 -8723 1484 -8689
rect -1546 -9758 -1512 -8782
rect 1512 -9758 1546 -8782
rect -1484 -9851 1484 -9817
rect -1484 -9959 1484 -9925
rect -1546 -10994 -1512 -10018
rect 1512 -10994 1546 -10018
rect -1484 -11087 1484 -11053
rect -1484 -11195 1484 -11161
rect -1546 -12230 -1512 -11254
rect 1512 -12230 1546 -11254
rect -1484 -12323 1484 -12289
rect -1484 -12431 1484 -12397
rect -1546 -13466 -1512 -12490
rect 1512 -13466 1546 -12490
rect -1484 -13559 1484 -13525
rect -1484 -13667 1484 -13633
rect -1546 -14702 -1512 -13726
rect 1512 -14702 1546 -13726
rect -1484 -14795 1484 -14761
rect -1484 -14903 1484 -14869
rect -1546 -15938 -1512 -14962
rect 1512 -15938 1546 -14962
rect -1484 -16031 1484 -15997
rect -1484 -16139 1484 -16105
rect -1546 -17174 -1512 -16198
rect 1512 -17174 1546 -16198
rect -1484 -17267 1484 -17233
rect -1484 -17375 1484 -17341
rect -1546 -18410 -1512 -17434
rect 1512 -18410 1546 -17434
rect -1484 -18503 1484 -18469
rect -1484 -18611 1484 -18577
rect -1546 -19646 -1512 -18670
rect 1512 -19646 1546 -18670
rect -1484 -19739 1484 -19705
rect -1484 -19847 1484 -19813
rect -1546 -20882 -1512 -19906
rect 1512 -20882 1546 -19906
rect -1484 -20975 1484 -20941
rect -1484 -21083 1484 -21049
rect -1546 -22118 -1512 -21142
rect 1512 -22118 1546 -21142
rect -1484 -22211 1484 -22177
rect -1484 -22319 1484 -22285
rect -1546 -23354 -1512 -22378
rect 1512 -23354 1546 -22378
rect -1484 -23447 1484 -23413
rect -1484 -23555 1484 -23521
rect -1546 -24590 -1512 -23614
rect 1512 -24590 1546 -23614
rect -1484 -24683 1484 -24649
rect -1484 -24791 1484 -24757
rect -1546 -25826 -1512 -24850
rect 1512 -25826 1546 -24850
rect -1484 -25919 1484 -25885
rect -1484 -26027 1484 -25993
rect -1546 -27062 -1512 -26086
rect 1512 -27062 1546 -26086
rect -1484 -27155 1484 -27121
rect -1484 -27263 1484 -27229
rect -1546 -28298 -1512 -27322
rect 1512 -28298 1546 -27322
rect -1484 -28391 1484 -28357
rect -1484 -28499 1484 -28465
rect -1546 -29534 -1512 -28558
rect 1512 -29534 1546 -28558
rect -1484 -29627 1484 -29593
rect -1484 -29735 1484 -29701
rect -1546 -30770 -1512 -29794
rect 1512 -30770 1546 -29794
rect -1484 -30863 1484 -30829
rect -1484 -30971 1484 -30937
rect -1546 -32006 -1512 -31030
rect 1512 -32006 1546 -31030
rect -1484 -32099 1484 -32065
rect -1484 -32207 1484 -32173
rect -1546 -33242 -1512 -32266
rect 1512 -33242 1546 -32266
rect -1484 -33335 1484 -33301
rect -1484 -33443 1484 -33409
rect -1546 -34478 -1512 -33502
rect 1512 -34478 1546 -33502
rect -1484 -34571 1484 -34537
rect -1484 -34679 1484 -34645
rect -1546 -35714 -1512 -34738
rect 1512 -35714 1546 -34738
rect -1484 -35807 1484 -35773
rect -1484 -35915 1484 -35881
rect -1546 -36950 -1512 -35974
rect 1512 -36950 1546 -35974
rect -1484 -37043 1484 -37009
rect -1484 -37151 1484 -37117
rect -1546 -38186 -1512 -37210
rect 1512 -38186 1546 -37210
rect -1484 -38279 1484 -38245
rect -1484 -38387 1484 -38353
rect -1546 -39422 -1512 -38446
rect 1512 -39422 1546 -38446
rect -1484 -39515 1484 -39481
rect -1484 -39623 1484 -39589
rect -1546 -40658 -1512 -39682
rect 1512 -40658 1546 -39682
rect -1484 -40751 1484 -40717
rect -1484 -40859 1484 -40825
rect -1546 -41894 -1512 -40918
rect 1512 -41894 1546 -40918
rect -1484 -41987 1484 -41953
rect -1484 -42095 1484 -42061
rect -1546 -43130 -1512 -42154
rect 1512 -43130 1546 -42154
rect -1484 -43223 1484 -43189
rect -1484 -43331 1484 -43297
rect -1546 -44366 -1512 -43390
rect 1512 -44366 1546 -43390
rect -1484 -44459 1484 -44425
rect -1484 -44567 1484 -44533
rect -1546 -45602 -1512 -44626
rect 1512 -45602 1546 -44626
rect -1484 -45695 1484 -45661
rect -1484 -45803 1484 -45769
rect -1546 -46838 -1512 -45862
rect 1512 -46838 1546 -45862
rect -1484 -46931 1484 -46897
rect -1484 -47039 1484 -47005
rect -1546 -48074 -1512 -47098
rect 1512 -48074 1546 -47098
rect -1484 -48167 1484 -48133
rect -1484 -48275 1484 -48241
rect -1546 -49310 -1512 -48334
rect 1512 -49310 1546 -48334
rect -1484 -49403 1484 -49369
rect -1484 -49511 1484 -49477
rect -1546 -50546 -1512 -49570
rect 1512 -50546 1546 -49570
rect -1484 -50639 1484 -50605
rect -1484 -50747 1484 -50713
rect -1546 -51782 -1512 -50806
rect 1512 -51782 1546 -50806
rect -1484 -51875 1484 -51841
rect -1484 -51983 1484 -51949
rect -1546 -53018 -1512 -52042
rect 1512 -53018 1546 -52042
rect -1484 -53111 1484 -53077
rect -1484 -53219 1484 -53185
rect -1546 -54254 -1512 -53278
rect 1512 -54254 1546 -53278
rect -1484 -54347 1484 -54313
rect -1484 -54455 1484 -54421
rect -1546 -55490 -1512 -54514
rect 1512 -55490 1546 -54514
rect -1484 -55583 1484 -55549
rect -1484 -55691 1484 -55657
rect -1546 -56726 -1512 -55750
rect 1512 -56726 1546 -55750
rect -1484 -56819 1484 -56785
rect -1484 -56927 1484 -56893
rect -1546 -57962 -1512 -56986
rect 1512 -57962 1546 -56986
rect -1484 -58055 1484 -58021
rect -1484 -58163 1484 -58129
rect -1546 -59198 -1512 -58222
rect 1512 -59198 1546 -58222
rect -1484 -59291 1484 -59257
rect -1484 -59399 1484 -59365
rect -1546 -60434 -1512 -59458
rect 1512 -60434 1546 -59458
rect -1484 -60527 1484 -60493
rect -1484 -60635 1484 -60601
rect -1546 -61670 -1512 -60694
rect 1512 -61670 1546 -60694
rect -1484 -61763 1484 -61729
rect -1484 -61871 1484 -61837
rect -1546 -62906 -1512 -61930
rect 1512 -62906 1546 -61930
rect -1484 -62999 1484 -62965
<< metal1 >>
rect -1496 62999 1496 63005
rect -1496 62965 -1484 62999
rect 1484 62965 1496 62999
rect -1496 62959 1496 62965
rect -1552 62906 -1506 62918
rect -1552 61930 -1546 62906
rect -1512 61930 -1506 62906
rect -1552 61918 -1506 61930
rect 1506 62906 1552 62918
rect 1506 61930 1512 62906
rect 1546 61930 1552 62906
rect 1506 61918 1552 61930
rect -1496 61871 1496 61877
rect -1496 61837 -1484 61871
rect 1484 61837 1496 61871
rect -1496 61831 1496 61837
rect -1496 61763 1496 61769
rect -1496 61729 -1484 61763
rect 1484 61729 1496 61763
rect -1496 61723 1496 61729
rect -1552 61670 -1506 61682
rect -1552 60694 -1546 61670
rect -1512 60694 -1506 61670
rect -1552 60682 -1506 60694
rect 1506 61670 1552 61682
rect 1506 60694 1512 61670
rect 1546 60694 1552 61670
rect 1506 60682 1552 60694
rect -1496 60635 1496 60641
rect -1496 60601 -1484 60635
rect 1484 60601 1496 60635
rect -1496 60595 1496 60601
rect -1496 60527 1496 60533
rect -1496 60493 -1484 60527
rect 1484 60493 1496 60527
rect -1496 60487 1496 60493
rect -1552 60434 -1506 60446
rect -1552 59458 -1546 60434
rect -1512 59458 -1506 60434
rect -1552 59446 -1506 59458
rect 1506 60434 1552 60446
rect 1506 59458 1512 60434
rect 1546 59458 1552 60434
rect 1506 59446 1552 59458
rect -1496 59399 1496 59405
rect -1496 59365 -1484 59399
rect 1484 59365 1496 59399
rect -1496 59359 1496 59365
rect -1496 59291 1496 59297
rect -1496 59257 -1484 59291
rect 1484 59257 1496 59291
rect -1496 59251 1496 59257
rect -1552 59198 -1506 59210
rect -1552 58222 -1546 59198
rect -1512 58222 -1506 59198
rect -1552 58210 -1506 58222
rect 1506 59198 1552 59210
rect 1506 58222 1512 59198
rect 1546 58222 1552 59198
rect 1506 58210 1552 58222
rect -1496 58163 1496 58169
rect -1496 58129 -1484 58163
rect 1484 58129 1496 58163
rect -1496 58123 1496 58129
rect -1496 58055 1496 58061
rect -1496 58021 -1484 58055
rect 1484 58021 1496 58055
rect -1496 58015 1496 58021
rect -1552 57962 -1506 57974
rect -1552 56986 -1546 57962
rect -1512 56986 -1506 57962
rect -1552 56974 -1506 56986
rect 1506 57962 1552 57974
rect 1506 56986 1512 57962
rect 1546 56986 1552 57962
rect 1506 56974 1552 56986
rect -1496 56927 1496 56933
rect -1496 56893 -1484 56927
rect 1484 56893 1496 56927
rect -1496 56887 1496 56893
rect -1496 56819 1496 56825
rect -1496 56785 -1484 56819
rect 1484 56785 1496 56819
rect -1496 56779 1496 56785
rect -1552 56726 -1506 56738
rect -1552 55750 -1546 56726
rect -1512 55750 -1506 56726
rect -1552 55738 -1506 55750
rect 1506 56726 1552 56738
rect 1506 55750 1512 56726
rect 1546 55750 1552 56726
rect 1506 55738 1552 55750
rect -1496 55691 1496 55697
rect -1496 55657 -1484 55691
rect 1484 55657 1496 55691
rect -1496 55651 1496 55657
rect -1496 55583 1496 55589
rect -1496 55549 -1484 55583
rect 1484 55549 1496 55583
rect -1496 55543 1496 55549
rect -1552 55490 -1506 55502
rect -1552 54514 -1546 55490
rect -1512 54514 -1506 55490
rect -1552 54502 -1506 54514
rect 1506 55490 1552 55502
rect 1506 54514 1512 55490
rect 1546 54514 1552 55490
rect 1506 54502 1552 54514
rect -1496 54455 1496 54461
rect -1496 54421 -1484 54455
rect 1484 54421 1496 54455
rect -1496 54415 1496 54421
rect -1496 54347 1496 54353
rect -1496 54313 -1484 54347
rect 1484 54313 1496 54347
rect -1496 54307 1496 54313
rect -1552 54254 -1506 54266
rect -1552 53278 -1546 54254
rect -1512 53278 -1506 54254
rect -1552 53266 -1506 53278
rect 1506 54254 1552 54266
rect 1506 53278 1512 54254
rect 1546 53278 1552 54254
rect 1506 53266 1552 53278
rect -1496 53219 1496 53225
rect -1496 53185 -1484 53219
rect 1484 53185 1496 53219
rect -1496 53179 1496 53185
rect -1496 53111 1496 53117
rect -1496 53077 -1484 53111
rect 1484 53077 1496 53111
rect -1496 53071 1496 53077
rect -1552 53018 -1506 53030
rect -1552 52042 -1546 53018
rect -1512 52042 -1506 53018
rect -1552 52030 -1506 52042
rect 1506 53018 1552 53030
rect 1506 52042 1512 53018
rect 1546 52042 1552 53018
rect 1506 52030 1552 52042
rect -1496 51983 1496 51989
rect -1496 51949 -1484 51983
rect 1484 51949 1496 51983
rect -1496 51943 1496 51949
rect -1496 51875 1496 51881
rect -1496 51841 -1484 51875
rect 1484 51841 1496 51875
rect -1496 51835 1496 51841
rect -1552 51782 -1506 51794
rect -1552 50806 -1546 51782
rect -1512 50806 -1506 51782
rect -1552 50794 -1506 50806
rect 1506 51782 1552 51794
rect 1506 50806 1512 51782
rect 1546 50806 1552 51782
rect 1506 50794 1552 50806
rect -1496 50747 1496 50753
rect -1496 50713 -1484 50747
rect 1484 50713 1496 50747
rect -1496 50707 1496 50713
rect -1496 50639 1496 50645
rect -1496 50605 -1484 50639
rect 1484 50605 1496 50639
rect -1496 50599 1496 50605
rect -1552 50546 -1506 50558
rect -1552 49570 -1546 50546
rect -1512 49570 -1506 50546
rect -1552 49558 -1506 49570
rect 1506 50546 1552 50558
rect 1506 49570 1512 50546
rect 1546 49570 1552 50546
rect 1506 49558 1552 49570
rect -1496 49511 1496 49517
rect -1496 49477 -1484 49511
rect 1484 49477 1496 49511
rect -1496 49471 1496 49477
rect -1496 49403 1496 49409
rect -1496 49369 -1484 49403
rect 1484 49369 1496 49403
rect -1496 49363 1496 49369
rect -1552 49310 -1506 49322
rect -1552 48334 -1546 49310
rect -1512 48334 -1506 49310
rect -1552 48322 -1506 48334
rect 1506 49310 1552 49322
rect 1506 48334 1512 49310
rect 1546 48334 1552 49310
rect 1506 48322 1552 48334
rect -1496 48275 1496 48281
rect -1496 48241 -1484 48275
rect 1484 48241 1496 48275
rect -1496 48235 1496 48241
rect -1496 48167 1496 48173
rect -1496 48133 -1484 48167
rect 1484 48133 1496 48167
rect -1496 48127 1496 48133
rect -1552 48074 -1506 48086
rect -1552 47098 -1546 48074
rect -1512 47098 -1506 48074
rect -1552 47086 -1506 47098
rect 1506 48074 1552 48086
rect 1506 47098 1512 48074
rect 1546 47098 1552 48074
rect 1506 47086 1552 47098
rect -1496 47039 1496 47045
rect -1496 47005 -1484 47039
rect 1484 47005 1496 47039
rect -1496 46999 1496 47005
rect -1496 46931 1496 46937
rect -1496 46897 -1484 46931
rect 1484 46897 1496 46931
rect -1496 46891 1496 46897
rect -1552 46838 -1506 46850
rect -1552 45862 -1546 46838
rect -1512 45862 -1506 46838
rect -1552 45850 -1506 45862
rect 1506 46838 1552 46850
rect 1506 45862 1512 46838
rect 1546 45862 1552 46838
rect 1506 45850 1552 45862
rect -1496 45803 1496 45809
rect -1496 45769 -1484 45803
rect 1484 45769 1496 45803
rect -1496 45763 1496 45769
rect -1496 45695 1496 45701
rect -1496 45661 -1484 45695
rect 1484 45661 1496 45695
rect -1496 45655 1496 45661
rect -1552 45602 -1506 45614
rect -1552 44626 -1546 45602
rect -1512 44626 -1506 45602
rect -1552 44614 -1506 44626
rect 1506 45602 1552 45614
rect 1506 44626 1512 45602
rect 1546 44626 1552 45602
rect 1506 44614 1552 44626
rect -1496 44567 1496 44573
rect -1496 44533 -1484 44567
rect 1484 44533 1496 44567
rect -1496 44527 1496 44533
rect -1496 44459 1496 44465
rect -1496 44425 -1484 44459
rect 1484 44425 1496 44459
rect -1496 44419 1496 44425
rect -1552 44366 -1506 44378
rect -1552 43390 -1546 44366
rect -1512 43390 -1506 44366
rect -1552 43378 -1506 43390
rect 1506 44366 1552 44378
rect 1506 43390 1512 44366
rect 1546 43390 1552 44366
rect 1506 43378 1552 43390
rect -1496 43331 1496 43337
rect -1496 43297 -1484 43331
rect 1484 43297 1496 43331
rect -1496 43291 1496 43297
rect -1496 43223 1496 43229
rect -1496 43189 -1484 43223
rect 1484 43189 1496 43223
rect -1496 43183 1496 43189
rect -1552 43130 -1506 43142
rect -1552 42154 -1546 43130
rect -1512 42154 -1506 43130
rect -1552 42142 -1506 42154
rect 1506 43130 1552 43142
rect 1506 42154 1512 43130
rect 1546 42154 1552 43130
rect 1506 42142 1552 42154
rect -1496 42095 1496 42101
rect -1496 42061 -1484 42095
rect 1484 42061 1496 42095
rect -1496 42055 1496 42061
rect -1496 41987 1496 41993
rect -1496 41953 -1484 41987
rect 1484 41953 1496 41987
rect -1496 41947 1496 41953
rect -1552 41894 -1506 41906
rect -1552 40918 -1546 41894
rect -1512 40918 -1506 41894
rect -1552 40906 -1506 40918
rect 1506 41894 1552 41906
rect 1506 40918 1512 41894
rect 1546 40918 1552 41894
rect 1506 40906 1552 40918
rect -1496 40859 1496 40865
rect -1496 40825 -1484 40859
rect 1484 40825 1496 40859
rect -1496 40819 1496 40825
rect -1496 40751 1496 40757
rect -1496 40717 -1484 40751
rect 1484 40717 1496 40751
rect -1496 40711 1496 40717
rect -1552 40658 -1506 40670
rect -1552 39682 -1546 40658
rect -1512 39682 -1506 40658
rect -1552 39670 -1506 39682
rect 1506 40658 1552 40670
rect 1506 39682 1512 40658
rect 1546 39682 1552 40658
rect 1506 39670 1552 39682
rect -1496 39623 1496 39629
rect -1496 39589 -1484 39623
rect 1484 39589 1496 39623
rect -1496 39583 1496 39589
rect -1496 39515 1496 39521
rect -1496 39481 -1484 39515
rect 1484 39481 1496 39515
rect -1496 39475 1496 39481
rect -1552 39422 -1506 39434
rect -1552 38446 -1546 39422
rect -1512 38446 -1506 39422
rect -1552 38434 -1506 38446
rect 1506 39422 1552 39434
rect 1506 38446 1512 39422
rect 1546 38446 1552 39422
rect 1506 38434 1552 38446
rect -1496 38387 1496 38393
rect -1496 38353 -1484 38387
rect 1484 38353 1496 38387
rect -1496 38347 1496 38353
rect -1496 38279 1496 38285
rect -1496 38245 -1484 38279
rect 1484 38245 1496 38279
rect -1496 38239 1496 38245
rect -1552 38186 -1506 38198
rect -1552 37210 -1546 38186
rect -1512 37210 -1506 38186
rect -1552 37198 -1506 37210
rect 1506 38186 1552 38198
rect 1506 37210 1512 38186
rect 1546 37210 1552 38186
rect 1506 37198 1552 37210
rect -1496 37151 1496 37157
rect -1496 37117 -1484 37151
rect 1484 37117 1496 37151
rect -1496 37111 1496 37117
rect -1496 37043 1496 37049
rect -1496 37009 -1484 37043
rect 1484 37009 1496 37043
rect -1496 37003 1496 37009
rect -1552 36950 -1506 36962
rect -1552 35974 -1546 36950
rect -1512 35974 -1506 36950
rect -1552 35962 -1506 35974
rect 1506 36950 1552 36962
rect 1506 35974 1512 36950
rect 1546 35974 1552 36950
rect 1506 35962 1552 35974
rect -1496 35915 1496 35921
rect -1496 35881 -1484 35915
rect 1484 35881 1496 35915
rect -1496 35875 1496 35881
rect -1496 35807 1496 35813
rect -1496 35773 -1484 35807
rect 1484 35773 1496 35807
rect -1496 35767 1496 35773
rect -1552 35714 -1506 35726
rect -1552 34738 -1546 35714
rect -1512 34738 -1506 35714
rect -1552 34726 -1506 34738
rect 1506 35714 1552 35726
rect 1506 34738 1512 35714
rect 1546 34738 1552 35714
rect 1506 34726 1552 34738
rect -1496 34679 1496 34685
rect -1496 34645 -1484 34679
rect 1484 34645 1496 34679
rect -1496 34639 1496 34645
rect -1496 34571 1496 34577
rect -1496 34537 -1484 34571
rect 1484 34537 1496 34571
rect -1496 34531 1496 34537
rect -1552 34478 -1506 34490
rect -1552 33502 -1546 34478
rect -1512 33502 -1506 34478
rect -1552 33490 -1506 33502
rect 1506 34478 1552 34490
rect 1506 33502 1512 34478
rect 1546 33502 1552 34478
rect 1506 33490 1552 33502
rect -1496 33443 1496 33449
rect -1496 33409 -1484 33443
rect 1484 33409 1496 33443
rect -1496 33403 1496 33409
rect -1496 33335 1496 33341
rect -1496 33301 -1484 33335
rect 1484 33301 1496 33335
rect -1496 33295 1496 33301
rect -1552 33242 -1506 33254
rect -1552 32266 -1546 33242
rect -1512 32266 -1506 33242
rect -1552 32254 -1506 32266
rect 1506 33242 1552 33254
rect 1506 32266 1512 33242
rect 1546 32266 1552 33242
rect 1506 32254 1552 32266
rect -1496 32207 1496 32213
rect -1496 32173 -1484 32207
rect 1484 32173 1496 32207
rect -1496 32167 1496 32173
rect -1496 32099 1496 32105
rect -1496 32065 -1484 32099
rect 1484 32065 1496 32099
rect -1496 32059 1496 32065
rect -1552 32006 -1506 32018
rect -1552 31030 -1546 32006
rect -1512 31030 -1506 32006
rect -1552 31018 -1506 31030
rect 1506 32006 1552 32018
rect 1506 31030 1512 32006
rect 1546 31030 1552 32006
rect 1506 31018 1552 31030
rect -1496 30971 1496 30977
rect -1496 30937 -1484 30971
rect 1484 30937 1496 30971
rect -1496 30931 1496 30937
rect -1496 30863 1496 30869
rect -1496 30829 -1484 30863
rect 1484 30829 1496 30863
rect -1496 30823 1496 30829
rect -1552 30770 -1506 30782
rect -1552 29794 -1546 30770
rect -1512 29794 -1506 30770
rect -1552 29782 -1506 29794
rect 1506 30770 1552 30782
rect 1506 29794 1512 30770
rect 1546 29794 1552 30770
rect 1506 29782 1552 29794
rect -1496 29735 1496 29741
rect -1496 29701 -1484 29735
rect 1484 29701 1496 29735
rect -1496 29695 1496 29701
rect -1496 29627 1496 29633
rect -1496 29593 -1484 29627
rect 1484 29593 1496 29627
rect -1496 29587 1496 29593
rect -1552 29534 -1506 29546
rect -1552 28558 -1546 29534
rect -1512 28558 -1506 29534
rect -1552 28546 -1506 28558
rect 1506 29534 1552 29546
rect 1506 28558 1512 29534
rect 1546 28558 1552 29534
rect 1506 28546 1552 28558
rect -1496 28499 1496 28505
rect -1496 28465 -1484 28499
rect 1484 28465 1496 28499
rect -1496 28459 1496 28465
rect -1496 28391 1496 28397
rect -1496 28357 -1484 28391
rect 1484 28357 1496 28391
rect -1496 28351 1496 28357
rect -1552 28298 -1506 28310
rect -1552 27322 -1546 28298
rect -1512 27322 -1506 28298
rect -1552 27310 -1506 27322
rect 1506 28298 1552 28310
rect 1506 27322 1512 28298
rect 1546 27322 1552 28298
rect 1506 27310 1552 27322
rect -1496 27263 1496 27269
rect -1496 27229 -1484 27263
rect 1484 27229 1496 27263
rect -1496 27223 1496 27229
rect -1496 27155 1496 27161
rect -1496 27121 -1484 27155
rect 1484 27121 1496 27155
rect -1496 27115 1496 27121
rect -1552 27062 -1506 27074
rect -1552 26086 -1546 27062
rect -1512 26086 -1506 27062
rect -1552 26074 -1506 26086
rect 1506 27062 1552 27074
rect 1506 26086 1512 27062
rect 1546 26086 1552 27062
rect 1506 26074 1552 26086
rect -1496 26027 1496 26033
rect -1496 25993 -1484 26027
rect 1484 25993 1496 26027
rect -1496 25987 1496 25993
rect -1496 25919 1496 25925
rect -1496 25885 -1484 25919
rect 1484 25885 1496 25919
rect -1496 25879 1496 25885
rect -1552 25826 -1506 25838
rect -1552 24850 -1546 25826
rect -1512 24850 -1506 25826
rect -1552 24838 -1506 24850
rect 1506 25826 1552 25838
rect 1506 24850 1512 25826
rect 1546 24850 1552 25826
rect 1506 24838 1552 24850
rect -1496 24791 1496 24797
rect -1496 24757 -1484 24791
rect 1484 24757 1496 24791
rect -1496 24751 1496 24757
rect -1496 24683 1496 24689
rect -1496 24649 -1484 24683
rect 1484 24649 1496 24683
rect -1496 24643 1496 24649
rect -1552 24590 -1506 24602
rect -1552 23614 -1546 24590
rect -1512 23614 -1506 24590
rect -1552 23602 -1506 23614
rect 1506 24590 1552 24602
rect 1506 23614 1512 24590
rect 1546 23614 1552 24590
rect 1506 23602 1552 23614
rect -1496 23555 1496 23561
rect -1496 23521 -1484 23555
rect 1484 23521 1496 23555
rect -1496 23515 1496 23521
rect -1496 23447 1496 23453
rect -1496 23413 -1484 23447
rect 1484 23413 1496 23447
rect -1496 23407 1496 23413
rect -1552 23354 -1506 23366
rect -1552 22378 -1546 23354
rect -1512 22378 -1506 23354
rect -1552 22366 -1506 22378
rect 1506 23354 1552 23366
rect 1506 22378 1512 23354
rect 1546 22378 1552 23354
rect 1506 22366 1552 22378
rect -1496 22319 1496 22325
rect -1496 22285 -1484 22319
rect 1484 22285 1496 22319
rect -1496 22279 1496 22285
rect -1496 22211 1496 22217
rect -1496 22177 -1484 22211
rect 1484 22177 1496 22211
rect -1496 22171 1496 22177
rect -1552 22118 -1506 22130
rect -1552 21142 -1546 22118
rect -1512 21142 -1506 22118
rect -1552 21130 -1506 21142
rect 1506 22118 1552 22130
rect 1506 21142 1512 22118
rect 1546 21142 1552 22118
rect 1506 21130 1552 21142
rect -1496 21083 1496 21089
rect -1496 21049 -1484 21083
rect 1484 21049 1496 21083
rect -1496 21043 1496 21049
rect -1496 20975 1496 20981
rect -1496 20941 -1484 20975
rect 1484 20941 1496 20975
rect -1496 20935 1496 20941
rect -1552 20882 -1506 20894
rect -1552 19906 -1546 20882
rect -1512 19906 -1506 20882
rect -1552 19894 -1506 19906
rect 1506 20882 1552 20894
rect 1506 19906 1512 20882
rect 1546 19906 1552 20882
rect 1506 19894 1552 19906
rect -1496 19847 1496 19853
rect -1496 19813 -1484 19847
rect 1484 19813 1496 19847
rect -1496 19807 1496 19813
rect -1496 19739 1496 19745
rect -1496 19705 -1484 19739
rect 1484 19705 1496 19739
rect -1496 19699 1496 19705
rect -1552 19646 -1506 19658
rect -1552 18670 -1546 19646
rect -1512 18670 -1506 19646
rect -1552 18658 -1506 18670
rect 1506 19646 1552 19658
rect 1506 18670 1512 19646
rect 1546 18670 1552 19646
rect 1506 18658 1552 18670
rect -1496 18611 1496 18617
rect -1496 18577 -1484 18611
rect 1484 18577 1496 18611
rect -1496 18571 1496 18577
rect -1496 18503 1496 18509
rect -1496 18469 -1484 18503
rect 1484 18469 1496 18503
rect -1496 18463 1496 18469
rect -1552 18410 -1506 18422
rect -1552 17434 -1546 18410
rect -1512 17434 -1506 18410
rect -1552 17422 -1506 17434
rect 1506 18410 1552 18422
rect 1506 17434 1512 18410
rect 1546 17434 1552 18410
rect 1506 17422 1552 17434
rect -1496 17375 1496 17381
rect -1496 17341 -1484 17375
rect 1484 17341 1496 17375
rect -1496 17335 1496 17341
rect -1496 17267 1496 17273
rect -1496 17233 -1484 17267
rect 1484 17233 1496 17267
rect -1496 17227 1496 17233
rect -1552 17174 -1506 17186
rect -1552 16198 -1546 17174
rect -1512 16198 -1506 17174
rect -1552 16186 -1506 16198
rect 1506 17174 1552 17186
rect 1506 16198 1512 17174
rect 1546 16198 1552 17174
rect 1506 16186 1552 16198
rect -1496 16139 1496 16145
rect -1496 16105 -1484 16139
rect 1484 16105 1496 16139
rect -1496 16099 1496 16105
rect -1496 16031 1496 16037
rect -1496 15997 -1484 16031
rect 1484 15997 1496 16031
rect -1496 15991 1496 15997
rect -1552 15938 -1506 15950
rect -1552 14962 -1546 15938
rect -1512 14962 -1506 15938
rect -1552 14950 -1506 14962
rect 1506 15938 1552 15950
rect 1506 14962 1512 15938
rect 1546 14962 1552 15938
rect 1506 14950 1552 14962
rect -1496 14903 1496 14909
rect -1496 14869 -1484 14903
rect 1484 14869 1496 14903
rect -1496 14863 1496 14869
rect -1496 14795 1496 14801
rect -1496 14761 -1484 14795
rect 1484 14761 1496 14795
rect -1496 14755 1496 14761
rect -1552 14702 -1506 14714
rect -1552 13726 -1546 14702
rect -1512 13726 -1506 14702
rect -1552 13714 -1506 13726
rect 1506 14702 1552 14714
rect 1506 13726 1512 14702
rect 1546 13726 1552 14702
rect 1506 13714 1552 13726
rect -1496 13667 1496 13673
rect -1496 13633 -1484 13667
rect 1484 13633 1496 13667
rect -1496 13627 1496 13633
rect -1496 13559 1496 13565
rect -1496 13525 -1484 13559
rect 1484 13525 1496 13559
rect -1496 13519 1496 13525
rect -1552 13466 -1506 13478
rect -1552 12490 -1546 13466
rect -1512 12490 -1506 13466
rect -1552 12478 -1506 12490
rect 1506 13466 1552 13478
rect 1506 12490 1512 13466
rect 1546 12490 1552 13466
rect 1506 12478 1552 12490
rect -1496 12431 1496 12437
rect -1496 12397 -1484 12431
rect 1484 12397 1496 12431
rect -1496 12391 1496 12397
rect -1496 12323 1496 12329
rect -1496 12289 -1484 12323
rect 1484 12289 1496 12323
rect -1496 12283 1496 12289
rect -1552 12230 -1506 12242
rect -1552 11254 -1546 12230
rect -1512 11254 -1506 12230
rect -1552 11242 -1506 11254
rect 1506 12230 1552 12242
rect 1506 11254 1512 12230
rect 1546 11254 1552 12230
rect 1506 11242 1552 11254
rect -1496 11195 1496 11201
rect -1496 11161 -1484 11195
rect 1484 11161 1496 11195
rect -1496 11155 1496 11161
rect -1496 11087 1496 11093
rect -1496 11053 -1484 11087
rect 1484 11053 1496 11087
rect -1496 11047 1496 11053
rect -1552 10994 -1506 11006
rect -1552 10018 -1546 10994
rect -1512 10018 -1506 10994
rect -1552 10006 -1506 10018
rect 1506 10994 1552 11006
rect 1506 10018 1512 10994
rect 1546 10018 1552 10994
rect 1506 10006 1552 10018
rect -1496 9959 1496 9965
rect -1496 9925 -1484 9959
rect 1484 9925 1496 9959
rect -1496 9919 1496 9925
rect -1496 9851 1496 9857
rect -1496 9817 -1484 9851
rect 1484 9817 1496 9851
rect -1496 9811 1496 9817
rect -1552 9758 -1506 9770
rect -1552 8782 -1546 9758
rect -1512 8782 -1506 9758
rect -1552 8770 -1506 8782
rect 1506 9758 1552 9770
rect 1506 8782 1512 9758
rect 1546 8782 1552 9758
rect 1506 8770 1552 8782
rect -1496 8723 1496 8729
rect -1496 8689 -1484 8723
rect 1484 8689 1496 8723
rect -1496 8683 1496 8689
rect -1496 8615 1496 8621
rect -1496 8581 -1484 8615
rect 1484 8581 1496 8615
rect -1496 8575 1496 8581
rect -1552 8522 -1506 8534
rect -1552 7546 -1546 8522
rect -1512 7546 -1506 8522
rect -1552 7534 -1506 7546
rect 1506 8522 1552 8534
rect 1506 7546 1512 8522
rect 1546 7546 1552 8522
rect 1506 7534 1552 7546
rect -1496 7487 1496 7493
rect -1496 7453 -1484 7487
rect 1484 7453 1496 7487
rect -1496 7447 1496 7453
rect -1496 7379 1496 7385
rect -1496 7345 -1484 7379
rect 1484 7345 1496 7379
rect -1496 7339 1496 7345
rect -1552 7286 -1506 7298
rect -1552 6310 -1546 7286
rect -1512 6310 -1506 7286
rect -1552 6298 -1506 6310
rect 1506 7286 1552 7298
rect 1506 6310 1512 7286
rect 1546 6310 1552 7286
rect 1506 6298 1552 6310
rect -1496 6251 1496 6257
rect -1496 6217 -1484 6251
rect 1484 6217 1496 6251
rect -1496 6211 1496 6217
rect -1496 6143 1496 6149
rect -1496 6109 -1484 6143
rect 1484 6109 1496 6143
rect -1496 6103 1496 6109
rect -1552 6050 -1506 6062
rect -1552 5074 -1546 6050
rect -1512 5074 -1506 6050
rect -1552 5062 -1506 5074
rect 1506 6050 1552 6062
rect 1506 5074 1512 6050
rect 1546 5074 1552 6050
rect 1506 5062 1552 5074
rect -1496 5015 1496 5021
rect -1496 4981 -1484 5015
rect 1484 4981 1496 5015
rect -1496 4975 1496 4981
rect -1496 4907 1496 4913
rect -1496 4873 -1484 4907
rect 1484 4873 1496 4907
rect -1496 4867 1496 4873
rect -1552 4814 -1506 4826
rect -1552 3838 -1546 4814
rect -1512 3838 -1506 4814
rect -1552 3826 -1506 3838
rect 1506 4814 1552 4826
rect 1506 3838 1512 4814
rect 1546 3838 1552 4814
rect 1506 3826 1552 3838
rect -1496 3779 1496 3785
rect -1496 3745 -1484 3779
rect 1484 3745 1496 3779
rect -1496 3739 1496 3745
rect -1496 3671 1496 3677
rect -1496 3637 -1484 3671
rect 1484 3637 1496 3671
rect -1496 3631 1496 3637
rect -1552 3578 -1506 3590
rect -1552 2602 -1546 3578
rect -1512 2602 -1506 3578
rect -1552 2590 -1506 2602
rect 1506 3578 1552 3590
rect 1506 2602 1512 3578
rect 1546 2602 1552 3578
rect 1506 2590 1552 2602
rect -1496 2543 1496 2549
rect -1496 2509 -1484 2543
rect 1484 2509 1496 2543
rect -1496 2503 1496 2509
rect -1496 2435 1496 2441
rect -1496 2401 -1484 2435
rect 1484 2401 1496 2435
rect -1496 2395 1496 2401
rect -1552 2342 -1506 2354
rect -1552 1366 -1546 2342
rect -1512 1366 -1506 2342
rect -1552 1354 -1506 1366
rect 1506 2342 1552 2354
rect 1506 1366 1512 2342
rect 1546 1366 1552 2342
rect 1506 1354 1552 1366
rect -1496 1307 1496 1313
rect -1496 1273 -1484 1307
rect 1484 1273 1496 1307
rect -1496 1267 1496 1273
rect -1496 1199 1496 1205
rect -1496 1165 -1484 1199
rect 1484 1165 1496 1199
rect -1496 1159 1496 1165
rect -1552 1106 -1506 1118
rect -1552 130 -1546 1106
rect -1512 130 -1506 1106
rect -1552 118 -1506 130
rect 1506 1106 1552 1118
rect 1506 130 1512 1106
rect 1546 130 1552 1106
rect 1506 118 1552 130
rect -1496 71 1496 77
rect -1496 37 -1484 71
rect 1484 37 1496 71
rect -1496 31 1496 37
rect -1496 -37 1496 -31
rect -1496 -71 -1484 -37
rect 1484 -71 1496 -37
rect -1496 -77 1496 -71
rect -1552 -130 -1506 -118
rect -1552 -1106 -1546 -130
rect -1512 -1106 -1506 -130
rect -1552 -1118 -1506 -1106
rect 1506 -130 1552 -118
rect 1506 -1106 1512 -130
rect 1546 -1106 1552 -130
rect 1506 -1118 1552 -1106
rect -1496 -1165 1496 -1159
rect -1496 -1199 -1484 -1165
rect 1484 -1199 1496 -1165
rect -1496 -1205 1496 -1199
rect -1496 -1273 1496 -1267
rect -1496 -1307 -1484 -1273
rect 1484 -1307 1496 -1273
rect -1496 -1313 1496 -1307
rect -1552 -1366 -1506 -1354
rect -1552 -2342 -1546 -1366
rect -1512 -2342 -1506 -1366
rect -1552 -2354 -1506 -2342
rect 1506 -1366 1552 -1354
rect 1506 -2342 1512 -1366
rect 1546 -2342 1552 -1366
rect 1506 -2354 1552 -2342
rect -1496 -2401 1496 -2395
rect -1496 -2435 -1484 -2401
rect 1484 -2435 1496 -2401
rect -1496 -2441 1496 -2435
rect -1496 -2509 1496 -2503
rect -1496 -2543 -1484 -2509
rect 1484 -2543 1496 -2509
rect -1496 -2549 1496 -2543
rect -1552 -2602 -1506 -2590
rect -1552 -3578 -1546 -2602
rect -1512 -3578 -1506 -2602
rect -1552 -3590 -1506 -3578
rect 1506 -2602 1552 -2590
rect 1506 -3578 1512 -2602
rect 1546 -3578 1552 -2602
rect 1506 -3590 1552 -3578
rect -1496 -3637 1496 -3631
rect -1496 -3671 -1484 -3637
rect 1484 -3671 1496 -3637
rect -1496 -3677 1496 -3671
rect -1496 -3745 1496 -3739
rect -1496 -3779 -1484 -3745
rect 1484 -3779 1496 -3745
rect -1496 -3785 1496 -3779
rect -1552 -3838 -1506 -3826
rect -1552 -4814 -1546 -3838
rect -1512 -4814 -1506 -3838
rect -1552 -4826 -1506 -4814
rect 1506 -3838 1552 -3826
rect 1506 -4814 1512 -3838
rect 1546 -4814 1552 -3838
rect 1506 -4826 1552 -4814
rect -1496 -4873 1496 -4867
rect -1496 -4907 -1484 -4873
rect 1484 -4907 1496 -4873
rect -1496 -4913 1496 -4907
rect -1496 -4981 1496 -4975
rect -1496 -5015 -1484 -4981
rect 1484 -5015 1496 -4981
rect -1496 -5021 1496 -5015
rect -1552 -5074 -1506 -5062
rect -1552 -6050 -1546 -5074
rect -1512 -6050 -1506 -5074
rect -1552 -6062 -1506 -6050
rect 1506 -5074 1552 -5062
rect 1506 -6050 1512 -5074
rect 1546 -6050 1552 -5074
rect 1506 -6062 1552 -6050
rect -1496 -6109 1496 -6103
rect -1496 -6143 -1484 -6109
rect 1484 -6143 1496 -6109
rect -1496 -6149 1496 -6143
rect -1496 -6217 1496 -6211
rect -1496 -6251 -1484 -6217
rect 1484 -6251 1496 -6217
rect -1496 -6257 1496 -6251
rect -1552 -6310 -1506 -6298
rect -1552 -7286 -1546 -6310
rect -1512 -7286 -1506 -6310
rect -1552 -7298 -1506 -7286
rect 1506 -6310 1552 -6298
rect 1506 -7286 1512 -6310
rect 1546 -7286 1552 -6310
rect 1506 -7298 1552 -7286
rect -1496 -7345 1496 -7339
rect -1496 -7379 -1484 -7345
rect 1484 -7379 1496 -7345
rect -1496 -7385 1496 -7379
rect -1496 -7453 1496 -7447
rect -1496 -7487 -1484 -7453
rect 1484 -7487 1496 -7453
rect -1496 -7493 1496 -7487
rect -1552 -7546 -1506 -7534
rect -1552 -8522 -1546 -7546
rect -1512 -8522 -1506 -7546
rect -1552 -8534 -1506 -8522
rect 1506 -7546 1552 -7534
rect 1506 -8522 1512 -7546
rect 1546 -8522 1552 -7546
rect 1506 -8534 1552 -8522
rect -1496 -8581 1496 -8575
rect -1496 -8615 -1484 -8581
rect 1484 -8615 1496 -8581
rect -1496 -8621 1496 -8615
rect -1496 -8689 1496 -8683
rect -1496 -8723 -1484 -8689
rect 1484 -8723 1496 -8689
rect -1496 -8729 1496 -8723
rect -1552 -8782 -1506 -8770
rect -1552 -9758 -1546 -8782
rect -1512 -9758 -1506 -8782
rect -1552 -9770 -1506 -9758
rect 1506 -8782 1552 -8770
rect 1506 -9758 1512 -8782
rect 1546 -9758 1552 -8782
rect 1506 -9770 1552 -9758
rect -1496 -9817 1496 -9811
rect -1496 -9851 -1484 -9817
rect 1484 -9851 1496 -9817
rect -1496 -9857 1496 -9851
rect -1496 -9925 1496 -9919
rect -1496 -9959 -1484 -9925
rect 1484 -9959 1496 -9925
rect -1496 -9965 1496 -9959
rect -1552 -10018 -1506 -10006
rect -1552 -10994 -1546 -10018
rect -1512 -10994 -1506 -10018
rect -1552 -11006 -1506 -10994
rect 1506 -10018 1552 -10006
rect 1506 -10994 1512 -10018
rect 1546 -10994 1552 -10018
rect 1506 -11006 1552 -10994
rect -1496 -11053 1496 -11047
rect -1496 -11087 -1484 -11053
rect 1484 -11087 1496 -11053
rect -1496 -11093 1496 -11087
rect -1496 -11161 1496 -11155
rect -1496 -11195 -1484 -11161
rect 1484 -11195 1496 -11161
rect -1496 -11201 1496 -11195
rect -1552 -11254 -1506 -11242
rect -1552 -12230 -1546 -11254
rect -1512 -12230 -1506 -11254
rect -1552 -12242 -1506 -12230
rect 1506 -11254 1552 -11242
rect 1506 -12230 1512 -11254
rect 1546 -12230 1552 -11254
rect 1506 -12242 1552 -12230
rect -1496 -12289 1496 -12283
rect -1496 -12323 -1484 -12289
rect 1484 -12323 1496 -12289
rect -1496 -12329 1496 -12323
rect -1496 -12397 1496 -12391
rect -1496 -12431 -1484 -12397
rect 1484 -12431 1496 -12397
rect -1496 -12437 1496 -12431
rect -1552 -12490 -1506 -12478
rect -1552 -13466 -1546 -12490
rect -1512 -13466 -1506 -12490
rect -1552 -13478 -1506 -13466
rect 1506 -12490 1552 -12478
rect 1506 -13466 1512 -12490
rect 1546 -13466 1552 -12490
rect 1506 -13478 1552 -13466
rect -1496 -13525 1496 -13519
rect -1496 -13559 -1484 -13525
rect 1484 -13559 1496 -13525
rect -1496 -13565 1496 -13559
rect -1496 -13633 1496 -13627
rect -1496 -13667 -1484 -13633
rect 1484 -13667 1496 -13633
rect -1496 -13673 1496 -13667
rect -1552 -13726 -1506 -13714
rect -1552 -14702 -1546 -13726
rect -1512 -14702 -1506 -13726
rect -1552 -14714 -1506 -14702
rect 1506 -13726 1552 -13714
rect 1506 -14702 1512 -13726
rect 1546 -14702 1552 -13726
rect 1506 -14714 1552 -14702
rect -1496 -14761 1496 -14755
rect -1496 -14795 -1484 -14761
rect 1484 -14795 1496 -14761
rect -1496 -14801 1496 -14795
rect -1496 -14869 1496 -14863
rect -1496 -14903 -1484 -14869
rect 1484 -14903 1496 -14869
rect -1496 -14909 1496 -14903
rect -1552 -14962 -1506 -14950
rect -1552 -15938 -1546 -14962
rect -1512 -15938 -1506 -14962
rect -1552 -15950 -1506 -15938
rect 1506 -14962 1552 -14950
rect 1506 -15938 1512 -14962
rect 1546 -15938 1552 -14962
rect 1506 -15950 1552 -15938
rect -1496 -15997 1496 -15991
rect -1496 -16031 -1484 -15997
rect 1484 -16031 1496 -15997
rect -1496 -16037 1496 -16031
rect -1496 -16105 1496 -16099
rect -1496 -16139 -1484 -16105
rect 1484 -16139 1496 -16105
rect -1496 -16145 1496 -16139
rect -1552 -16198 -1506 -16186
rect -1552 -17174 -1546 -16198
rect -1512 -17174 -1506 -16198
rect -1552 -17186 -1506 -17174
rect 1506 -16198 1552 -16186
rect 1506 -17174 1512 -16198
rect 1546 -17174 1552 -16198
rect 1506 -17186 1552 -17174
rect -1496 -17233 1496 -17227
rect -1496 -17267 -1484 -17233
rect 1484 -17267 1496 -17233
rect -1496 -17273 1496 -17267
rect -1496 -17341 1496 -17335
rect -1496 -17375 -1484 -17341
rect 1484 -17375 1496 -17341
rect -1496 -17381 1496 -17375
rect -1552 -17434 -1506 -17422
rect -1552 -18410 -1546 -17434
rect -1512 -18410 -1506 -17434
rect -1552 -18422 -1506 -18410
rect 1506 -17434 1552 -17422
rect 1506 -18410 1512 -17434
rect 1546 -18410 1552 -17434
rect 1506 -18422 1552 -18410
rect -1496 -18469 1496 -18463
rect -1496 -18503 -1484 -18469
rect 1484 -18503 1496 -18469
rect -1496 -18509 1496 -18503
rect -1496 -18577 1496 -18571
rect -1496 -18611 -1484 -18577
rect 1484 -18611 1496 -18577
rect -1496 -18617 1496 -18611
rect -1552 -18670 -1506 -18658
rect -1552 -19646 -1546 -18670
rect -1512 -19646 -1506 -18670
rect -1552 -19658 -1506 -19646
rect 1506 -18670 1552 -18658
rect 1506 -19646 1512 -18670
rect 1546 -19646 1552 -18670
rect 1506 -19658 1552 -19646
rect -1496 -19705 1496 -19699
rect -1496 -19739 -1484 -19705
rect 1484 -19739 1496 -19705
rect -1496 -19745 1496 -19739
rect -1496 -19813 1496 -19807
rect -1496 -19847 -1484 -19813
rect 1484 -19847 1496 -19813
rect -1496 -19853 1496 -19847
rect -1552 -19906 -1506 -19894
rect -1552 -20882 -1546 -19906
rect -1512 -20882 -1506 -19906
rect -1552 -20894 -1506 -20882
rect 1506 -19906 1552 -19894
rect 1506 -20882 1512 -19906
rect 1546 -20882 1552 -19906
rect 1506 -20894 1552 -20882
rect -1496 -20941 1496 -20935
rect -1496 -20975 -1484 -20941
rect 1484 -20975 1496 -20941
rect -1496 -20981 1496 -20975
rect -1496 -21049 1496 -21043
rect -1496 -21083 -1484 -21049
rect 1484 -21083 1496 -21049
rect -1496 -21089 1496 -21083
rect -1552 -21142 -1506 -21130
rect -1552 -22118 -1546 -21142
rect -1512 -22118 -1506 -21142
rect -1552 -22130 -1506 -22118
rect 1506 -21142 1552 -21130
rect 1506 -22118 1512 -21142
rect 1546 -22118 1552 -21142
rect 1506 -22130 1552 -22118
rect -1496 -22177 1496 -22171
rect -1496 -22211 -1484 -22177
rect 1484 -22211 1496 -22177
rect -1496 -22217 1496 -22211
rect -1496 -22285 1496 -22279
rect -1496 -22319 -1484 -22285
rect 1484 -22319 1496 -22285
rect -1496 -22325 1496 -22319
rect -1552 -22378 -1506 -22366
rect -1552 -23354 -1546 -22378
rect -1512 -23354 -1506 -22378
rect -1552 -23366 -1506 -23354
rect 1506 -22378 1552 -22366
rect 1506 -23354 1512 -22378
rect 1546 -23354 1552 -22378
rect 1506 -23366 1552 -23354
rect -1496 -23413 1496 -23407
rect -1496 -23447 -1484 -23413
rect 1484 -23447 1496 -23413
rect -1496 -23453 1496 -23447
rect -1496 -23521 1496 -23515
rect -1496 -23555 -1484 -23521
rect 1484 -23555 1496 -23521
rect -1496 -23561 1496 -23555
rect -1552 -23614 -1506 -23602
rect -1552 -24590 -1546 -23614
rect -1512 -24590 -1506 -23614
rect -1552 -24602 -1506 -24590
rect 1506 -23614 1552 -23602
rect 1506 -24590 1512 -23614
rect 1546 -24590 1552 -23614
rect 1506 -24602 1552 -24590
rect -1496 -24649 1496 -24643
rect -1496 -24683 -1484 -24649
rect 1484 -24683 1496 -24649
rect -1496 -24689 1496 -24683
rect -1496 -24757 1496 -24751
rect -1496 -24791 -1484 -24757
rect 1484 -24791 1496 -24757
rect -1496 -24797 1496 -24791
rect -1552 -24850 -1506 -24838
rect -1552 -25826 -1546 -24850
rect -1512 -25826 -1506 -24850
rect -1552 -25838 -1506 -25826
rect 1506 -24850 1552 -24838
rect 1506 -25826 1512 -24850
rect 1546 -25826 1552 -24850
rect 1506 -25838 1552 -25826
rect -1496 -25885 1496 -25879
rect -1496 -25919 -1484 -25885
rect 1484 -25919 1496 -25885
rect -1496 -25925 1496 -25919
rect -1496 -25993 1496 -25987
rect -1496 -26027 -1484 -25993
rect 1484 -26027 1496 -25993
rect -1496 -26033 1496 -26027
rect -1552 -26086 -1506 -26074
rect -1552 -27062 -1546 -26086
rect -1512 -27062 -1506 -26086
rect -1552 -27074 -1506 -27062
rect 1506 -26086 1552 -26074
rect 1506 -27062 1512 -26086
rect 1546 -27062 1552 -26086
rect 1506 -27074 1552 -27062
rect -1496 -27121 1496 -27115
rect -1496 -27155 -1484 -27121
rect 1484 -27155 1496 -27121
rect -1496 -27161 1496 -27155
rect -1496 -27229 1496 -27223
rect -1496 -27263 -1484 -27229
rect 1484 -27263 1496 -27229
rect -1496 -27269 1496 -27263
rect -1552 -27322 -1506 -27310
rect -1552 -28298 -1546 -27322
rect -1512 -28298 -1506 -27322
rect -1552 -28310 -1506 -28298
rect 1506 -27322 1552 -27310
rect 1506 -28298 1512 -27322
rect 1546 -28298 1552 -27322
rect 1506 -28310 1552 -28298
rect -1496 -28357 1496 -28351
rect -1496 -28391 -1484 -28357
rect 1484 -28391 1496 -28357
rect -1496 -28397 1496 -28391
rect -1496 -28465 1496 -28459
rect -1496 -28499 -1484 -28465
rect 1484 -28499 1496 -28465
rect -1496 -28505 1496 -28499
rect -1552 -28558 -1506 -28546
rect -1552 -29534 -1546 -28558
rect -1512 -29534 -1506 -28558
rect -1552 -29546 -1506 -29534
rect 1506 -28558 1552 -28546
rect 1506 -29534 1512 -28558
rect 1546 -29534 1552 -28558
rect 1506 -29546 1552 -29534
rect -1496 -29593 1496 -29587
rect -1496 -29627 -1484 -29593
rect 1484 -29627 1496 -29593
rect -1496 -29633 1496 -29627
rect -1496 -29701 1496 -29695
rect -1496 -29735 -1484 -29701
rect 1484 -29735 1496 -29701
rect -1496 -29741 1496 -29735
rect -1552 -29794 -1506 -29782
rect -1552 -30770 -1546 -29794
rect -1512 -30770 -1506 -29794
rect -1552 -30782 -1506 -30770
rect 1506 -29794 1552 -29782
rect 1506 -30770 1512 -29794
rect 1546 -30770 1552 -29794
rect 1506 -30782 1552 -30770
rect -1496 -30829 1496 -30823
rect -1496 -30863 -1484 -30829
rect 1484 -30863 1496 -30829
rect -1496 -30869 1496 -30863
rect -1496 -30937 1496 -30931
rect -1496 -30971 -1484 -30937
rect 1484 -30971 1496 -30937
rect -1496 -30977 1496 -30971
rect -1552 -31030 -1506 -31018
rect -1552 -32006 -1546 -31030
rect -1512 -32006 -1506 -31030
rect -1552 -32018 -1506 -32006
rect 1506 -31030 1552 -31018
rect 1506 -32006 1512 -31030
rect 1546 -32006 1552 -31030
rect 1506 -32018 1552 -32006
rect -1496 -32065 1496 -32059
rect -1496 -32099 -1484 -32065
rect 1484 -32099 1496 -32065
rect -1496 -32105 1496 -32099
rect -1496 -32173 1496 -32167
rect -1496 -32207 -1484 -32173
rect 1484 -32207 1496 -32173
rect -1496 -32213 1496 -32207
rect -1552 -32266 -1506 -32254
rect -1552 -33242 -1546 -32266
rect -1512 -33242 -1506 -32266
rect -1552 -33254 -1506 -33242
rect 1506 -32266 1552 -32254
rect 1506 -33242 1512 -32266
rect 1546 -33242 1552 -32266
rect 1506 -33254 1552 -33242
rect -1496 -33301 1496 -33295
rect -1496 -33335 -1484 -33301
rect 1484 -33335 1496 -33301
rect -1496 -33341 1496 -33335
rect -1496 -33409 1496 -33403
rect -1496 -33443 -1484 -33409
rect 1484 -33443 1496 -33409
rect -1496 -33449 1496 -33443
rect -1552 -33502 -1506 -33490
rect -1552 -34478 -1546 -33502
rect -1512 -34478 -1506 -33502
rect -1552 -34490 -1506 -34478
rect 1506 -33502 1552 -33490
rect 1506 -34478 1512 -33502
rect 1546 -34478 1552 -33502
rect 1506 -34490 1552 -34478
rect -1496 -34537 1496 -34531
rect -1496 -34571 -1484 -34537
rect 1484 -34571 1496 -34537
rect -1496 -34577 1496 -34571
rect -1496 -34645 1496 -34639
rect -1496 -34679 -1484 -34645
rect 1484 -34679 1496 -34645
rect -1496 -34685 1496 -34679
rect -1552 -34738 -1506 -34726
rect -1552 -35714 -1546 -34738
rect -1512 -35714 -1506 -34738
rect -1552 -35726 -1506 -35714
rect 1506 -34738 1552 -34726
rect 1506 -35714 1512 -34738
rect 1546 -35714 1552 -34738
rect 1506 -35726 1552 -35714
rect -1496 -35773 1496 -35767
rect -1496 -35807 -1484 -35773
rect 1484 -35807 1496 -35773
rect -1496 -35813 1496 -35807
rect -1496 -35881 1496 -35875
rect -1496 -35915 -1484 -35881
rect 1484 -35915 1496 -35881
rect -1496 -35921 1496 -35915
rect -1552 -35974 -1506 -35962
rect -1552 -36950 -1546 -35974
rect -1512 -36950 -1506 -35974
rect -1552 -36962 -1506 -36950
rect 1506 -35974 1552 -35962
rect 1506 -36950 1512 -35974
rect 1546 -36950 1552 -35974
rect 1506 -36962 1552 -36950
rect -1496 -37009 1496 -37003
rect -1496 -37043 -1484 -37009
rect 1484 -37043 1496 -37009
rect -1496 -37049 1496 -37043
rect -1496 -37117 1496 -37111
rect -1496 -37151 -1484 -37117
rect 1484 -37151 1496 -37117
rect -1496 -37157 1496 -37151
rect -1552 -37210 -1506 -37198
rect -1552 -38186 -1546 -37210
rect -1512 -38186 -1506 -37210
rect -1552 -38198 -1506 -38186
rect 1506 -37210 1552 -37198
rect 1506 -38186 1512 -37210
rect 1546 -38186 1552 -37210
rect 1506 -38198 1552 -38186
rect -1496 -38245 1496 -38239
rect -1496 -38279 -1484 -38245
rect 1484 -38279 1496 -38245
rect -1496 -38285 1496 -38279
rect -1496 -38353 1496 -38347
rect -1496 -38387 -1484 -38353
rect 1484 -38387 1496 -38353
rect -1496 -38393 1496 -38387
rect -1552 -38446 -1506 -38434
rect -1552 -39422 -1546 -38446
rect -1512 -39422 -1506 -38446
rect -1552 -39434 -1506 -39422
rect 1506 -38446 1552 -38434
rect 1506 -39422 1512 -38446
rect 1546 -39422 1552 -38446
rect 1506 -39434 1552 -39422
rect -1496 -39481 1496 -39475
rect -1496 -39515 -1484 -39481
rect 1484 -39515 1496 -39481
rect -1496 -39521 1496 -39515
rect -1496 -39589 1496 -39583
rect -1496 -39623 -1484 -39589
rect 1484 -39623 1496 -39589
rect -1496 -39629 1496 -39623
rect -1552 -39682 -1506 -39670
rect -1552 -40658 -1546 -39682
rect -1512 -40658 -1506 -39682
rect -1552 -40670 -1506 -40658
rect 1506 -39682 1552 -39670
rect 1506 -40658 1512 -39682
rect 1546 -40658 1552 -39682
rect 1506 -40670 1552 -40658
rect -1496 -40717 1496 -40711
rect -1496 -40751 -1484 -40717
rect 1484 -40751 1496 -40717
rect -1496 -40757 1496 -40751
rect -1496 -40825 1496 -40819
rect -1496 -40859 -1484 -40825
rect 1484 -40859 1496 -40825
rect -1496 -40865 1496 -40859
rect -1552 -40918 -1506 -40906
rect -1552 -41894 -1546 -40918
rect -1512 -41894 -1506 -40918
rect -1552 -41906 -1506 -41894
rect 1506 -40918 1552 -40906
rect 1506 -41894 1512 -40918
rect 1546 -41894 1552 -40918
rect 1506 -41906 1552 -41894
rect -1496 -41953 1496 -41947
rect -1496 -41987 -1484 -41953
rect 1484 -41987 1496 -41953
rect -1496 -41993 1496 -41987
rect -1496 -42061 1496 -42055
rect -1496 -42095 -1484 -42061
rect 1484 -42095 1496 -42061
rect -1496 -42101 1496 -42095
rect -1552 -42154 -1506 -42142
rect -1552 -43130 -1546 -42154
rect -1512 -43130 -1506 -42154
rect -1552 -43142 -1506 -43130
rect 1506 -42154 1552 -42142
rect 1506 -43130 1512 -42154
rect 1546 -43130 1552 -42154
rect 1506 -43142 1552 -43130
rect -1496 -43189 1496 -43183
rect -1496 -43223 -1484 -43189
rect 1484 -43223 1496 -43189
rect -1496 -43229 1496 -43223
rect -1496 -43297 1496 -43291
rect -1496 -43331 -1484 -43297
rect 1484 -43331 1496 -43297
rect -1496 -43337 1496 -43331
rect -1552 -43390 -1506 -43378
rect -1552 -44366 -1546 -43390
rect -1512 -44366 -1506 -43390
rect -1552 -44378 -1506 -44366
rect 1506 -43390 1552 -43378
rect 1506 -44366 1512 -43390
rect 1546 -44366 1552 -43390
rect 1506 -44378 1552 -44366
rect -1496 -44425 1496 -44419
rect -1496 -44459 -1484 -44425
rect 1484 -44459 1496 -44425
rect -1496 -44465 1496 -44459
rect -1496 -44533 1496 -44527
rect -1496 -44567 -1484 -44533
rect 1484 -44567 1496 -44533
rect -1496 -44573 1496 -44567
rect -1552 -44626 -1506 -44614
rect -1552 -45602 -1546 -44626
rect -1512 -45602 -1506 -44626
rect -1552 -45614 -1506 -45602
rect 1506 -44626 1552 -44614
rect 1506 -45602 1512 -44626
rect 1546 -45602 1552 -44626
rect 1506 -45614 1552 -45602
rect -1496 -45661 1496 -45655
rect -1496 -45695 -1484 -45661
rect 1484 -45695 1496 -45661
rect -1496 -45701 1496 -45695
rect -1496 -45769 1496 -45763
rect -1496 -45803 -1484 -45769
rect 1484 -45803 1496 -45769
rect -1496 -45809 1496 -45803
rect -1552 -45862 -1506 -45850
rect -1552 -46838 -1546 -45862
rect -1512 -46838 -1506 -45862
rect -1552 -46850 -1506 -46838
rect 1506 -45862 1552 -45850
rect 1506 -46838 1512 -45862
rect 1546 -46838 1552 -45862
rect 1506 -46850 1552 -46838
rect -1496 -46897 1496 -46891
rect -1496 -46931 -1484 -46897
rect 1484 -46931 1496 -46897
rect -1496 -46937 1496 -46931
rect -1496 -47005 1496 -46999
rect -1496 -47039 -1484 -47005
rect 1484 -47039 1496 -47005
rect -1496 -47045 1496 -47039
rect -1552 -47098 -1506 -47086
rect -1552 -48074 -1546 -47098
rect -1512 -48074 -1506 -47098
rect -1552 -48086 -1506 -48074
rect 1506 -47098 1552 -47086
rect 1506 -48074 1512 -47098
rect 1546 -48074 1552 -47098
rect 1506 -48086 1552 -48074
rect -1496 -48133 1496 -48127
rect -1496 -48167 -1484 -48133
rect 1484 -48167 1496 -48133
rect -1496 -48173 1496 -48167
rect -1496 -48241 1496 -48235
rect -1496 -48275 -1484 -48241
rect 1484 -48275 1496 -48241
rect -1496 -48281 1496 -48275
rect -1552 -48334 -1506 -48322
rect -1552 -49310 -1546 -48334
rect -1512 -49310 -1506 -48334
rect -1552 -49322 -1506 -49310
rect 1506 -48334 1552 -48322
rect 1506 -49310 1512 -48334
rect 1546 -49310 1552 -48334
rect 1506 -49322 1552 -49310
rect -1496 -49369 1496 -49363
rect -1496 -49403 -1484 -49369
rect 1484 -49403 1496 -49369
rect -1496 -49409 1496 -49403
rect -1496 -49477 1496 -49471
rect -1496 -49511 -1484 -49477
rect 1484 -49511 1496 -49477
rect -1496 -49517 1496 -49511
rect -1552 -49570 -1506 -49558
rect -1552 -50546 -1546 -49570
rect -1512 -50546 -1506 -49570
rect -1552 -50558 -1506 -50546
rect 1506 -49570 1552 -49558
rect 1506 -50546 1512 -49570
rect 1546 -50546 1552 -49570
rect 1506 -50558 1552 -50546
rect -1496 -50605 1496 -50599
rect -1496 -50639 -1484 -50605
rect 1484 -50639 1496 -50605
rect -1496 -50645 1496 -50639
rect -1496 -50713 1496 -50707
rect -1496 -50747 -1484 -50713
rect 1484 -50747 1496 -50713
rect -1496 -50753 1496 -50747
rect -1552 -50806 -1506 -50794
rect -1552 -51782 -1546 -50806
rect -1512 -51782 -1506 -50806
rect -1552 -51794 -1506 -51782
rect 1506 -50806 1552 -50794
rect 1506 -51782 1512 -50806
rect 1546 -51782 1552 -50806
rect 1506 -51794 1552 -51782
rect -1496 -51841 1496 -51835
rect -1496 -51875 -1484 -51841
rect 1484 -51875 1496 -51841
rect -1496 -51881 1496 -51875
rect -1496 -51949 1496 -51943
rect -1496 -51983 -1484 -51949
rect 1484 -51983 1496 -51949
rect -1496 -51989 1496 -51983
rect -1552 -52042 -1506 -52030
rect -1552 -53018 -1546 -52042
rect -1512 -53018 -1506 -52042
rect -1552 -53030 -1506 -53018
rect 1506 -52042 1552 -52030
rect 1506 -53018 1512 -52042
rect 1546 -53018 1552 -52042
rect 1506 -53030 1552 -53018
rect -1496 -53077 1496 -53071
rect -1496 -53111 -1484 -53077
rect 1484 -53111 1496 -53077
rect -1496 -53117 1496 -53111
rect -1496 -53185 1496 -53179
rect -1496 -53219 -1484 -53185
rect 1484 -53219 1496 -53185
rect -1496 -53225 1496 -53219
rect -1552 -53278 -1506 -53266
rect -1552 -54254 -1546 -53278
rect -1512 -54254 -1506 -53278
rect -1552 -54266 -1506 -54254
rect 1506 -53278 1552 -53266
rect 1506 -54254 1512 -53278
rect 1546 -54254 1552 -53278
rect 1506 -54266 1552 -54254
rect -1496 -54313 1496 -54307
rect -1496 -54347 -1484 -54313
rect 1484 -54347 1496 -54313
rect -1496 -54353 1496 -54347
rect -1496 -54421 1496 -54415
rect -1496 -54455 -1484 -54421
rect 1484 -54455 1496 -54421
rect -1496 -54461 1496 -54455
rect -1552 -54514 -1506 -54502
rect -1552 -55490 -1546 -54514
rect -1512 -55490 -1506 -54514
rect -1552 -55502 -1506 -55490
rect 1506 -54514 1552 -54502
rect 1506 -55490 1512 -54514
rect 1546 -55490 1552 -54514
rect 1506 -55502 1552 -55490
rect -1496 -55549 1496 -55543
rect -1496 -55583 -1484 -55549
rect 1484 -55583 1496 -55549
rect -1496 -55589 1496 -55583
rect -1496 -55657 1496 -55651
rect -1496 -55691 -1484 -55657
rect 1484 -55691 1496 -55657
rect -1496 -55697 1496 -55691
rect -1552 -55750 -1506 -55738
rect -1552 -56726 -1546 -55750
rect -1512 -56726 -1506 -55750
rect -1552 -56738 -1506 -56726
rect 1506 -55750 1552 -55738
rect 1506 -56726 1512 -55750
rect 1546 -56726 1552 -55750
rect 1506 -56738 1552 -56726
rect -1496 -56785 1496 -56779
rect -1496 -56819 -1484 -56785
rect 1484 -56819 1496 -56785
rect -1496 -56825 1496 -56819
rect -1496 -56893 1496 -56887
rect -1496 -56927 -1484 -56893
rect 1484 -56927 1496 -56893
rect -1496 -56933 1496 -56927
rect -1552 -56986 -1506 -56974
rect -1552 -57962 -1546 -56986
rect -1512 -57962 -1506 -56986
rect -1552 -57974 -1506 -57962
rect 1506 -56986 1552 -56974
rect 1506 -57962 1512 -56986
rect 1546 -57962 1552 -56986
rect 1506 -57974 1552 -57962
rect -1496 -58021 1496 -58015
rect -1496 -58055 -1484 -58021
rect 1484 -58055 1496 -58021
rect -1496 -58061 1496 -58055
rect -1496 -58129 1496 -58123
rect -1496 -58163 -1484 -58129
rect 1484 -58163 1496 -58129
rect -1496 -58169 1496 -58163
rect -1552 -58222 -1506 -58210
rect -1552 -59198 -1546 -58222
rect -1512 -59198 -1506 -58222
rect -1552 -59210 -1506 -59198
rect 1506 -58222 1552 -58210
rect 1506 -59198 1512 -58222
rect 1546 -59198 1552 -58222
rect 1506 -59210 1552 -59198
rect -1496 -59257 1496 -59251
rect -1496 -59291 -1484 -59257
rect 1484 -59291 1496 -59257
rect -1496 -59297 1496 -59291
rect -1496 -59365 1496 -59359
rect -1496 -59399 -1484 -59365
rect 1484 -59399 1496 -59365
rect -1496 -59405 1496 -59399
rect -1552 -59458 -1506 -59446
rect -1552 -60434 -1546 -59458
rect -1512 -60434 -1506 -59458
rect -1552 -60446 -1506 -60434
rect 1506 -59458 1552 -59446
rect 1506 -60434 1512 -59458
rect 1546 -60434 1552 -59458
rect 1506 -60446 1552 -60434
rect -1496 -60493 1496 -60487
rect -1496 -60527 -1484 -60493
rect 1484 -60527 1496 -60493
rect -1496 -60533 1496 -60527
rect -1496 -60601 1496 -60595
rect -1496 -60635 -1484 -60601
rect 1484 -60635 1496 -60601
rect -1496 -60641 1496 -60635
rect -1552 -60694 -1506 -60682
rect -1552 -61670 -1546 -60694
rect -1512 -61670 -1506 -60694
rect -1552 -61682 -1506 -61670
rect 1506 -60694 1552 -60682
rect 1506 -61670 1512 -60694
rect 1546 -61670 1552 -60694
rect 1506 -61682 1552 -61670
rect -1496 -61729 1496 -61723
rect -1496 -61763 -1484 -61729
rect 1484 -61763 1496 -61729
rect -1496 -61769 1496 -61763
rect -1496 -61837 1496 -61831
rect -1496 -61871 -1484 -61837
rect 1484 -61871 1496 -61837
rect -1496 -61877 1496 -61871
rect -1552 -61930 -1506 -61918
rect -1552 -62906 -1546 -61930
rect -1512 -62906 -1506 -61930
rect -1552 -62918 -1506 -62906
rect 1506 -61930 1552 -61918
rect 1506 -62906 1512 -61930
rect 1546 -62906 1552 -61930
rect 1506 -62918 1552 -62906
rect -1496 -62965 1496 -62959
rect -1496 -62999 -1484 -62965
rect 1484 -62999 1496 -62965
rect -1496 -63005 1496 -62999
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 5.0 l 15.0 m 102 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
