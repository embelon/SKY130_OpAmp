* NGSPICE file created from opamp_cascode.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_SCE452 a_n158_n125# a_n100_n213# a_100_n125# VSUBS
X0 a_100_n125# a_n100_n213# a_n158_n125# VSUBS sky130_fd_pr__nfet_01v8 ad=0.363 pd=3.08 as=0.363 ps=3.08 w=1.25 l=1
**devattr s=14500,616 d=14500,616
C0 a_100_n125# a_n100_n213# 0.0322f
C1 a_n158_n125# a_n100_n213# 0.0322f
C2 a_n158_n125# a_100_n125# 0.0693f
C3 a_100_n125# VSUBS 0.151f
C4 a_n158_n125# VSUBS 0.151f
C5 a_n100_n213# VSUBS 0.664f
.ends

.subckt sky130_fd_pr__pfet_01v8_ZLZ7XS w_n1594_n600# a_n1500_n597# a_1500_n500# a_n1558_n500#
+ VSUBS
X0 a_1500_n500# a_n1500_n597# a_n1558_n500# w_n1594_n600# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
C0 a_n1558_n500# w_n1594_n600# 0.0187f
C1 a_n1500_n597# w_n1594_n600# 1.65f
C2 w_n1594_n600# a_1500_n500# 0.0187f
C3 a_n1500_n597# a_n1558_n500# 0.217f
C4 a_n1500_n597# a_1500_n500# 0.217f
C5 a_1500_n500# VSUBS 0.65f
C6 a_n1558_n500# VSUBS 0.65f
C7 a_n1500_n597# VSUBS 6.74f
C8 w_n1594_n600# VSUBS 11.5f
.ends

.subckt sky130_fd_pr__pfet_01v8_7DHACV w_n112_636# a_n33_n5541# a_n33_n8013# a_n76_736#
+ w_n112_1872# w_n112_4344# a_18_n500# a_18_n2972# a_18_n5444# a_n76_n1736# a_n33_3111#
+ a_n76_n4208# a_18_3208# a_n76_n7916# a_n33_n1833# a_18_6916# a_n76_5680# w_n112_n3072#
+ a_n33_n4305# a_n33_5583# a_n76_8152# w_n112_n6780# a_n33_8055# a_n33_n3069# a_n33_639#
+ w_n112_n9252# w_n112_3108# w_n112_6816# a_n33_n6777# a_n33_n597# a_n33_n9249# a_18_n1736#
+ a_18_n4208# a_18_n7916# a_n76_1972# a_n33_1875# w_n112_n600# a_n76_n6680# a_18_736#
+ a_n76_4444# a_18_5680# a_n33_4347# w_n112_n5544# a_n76_n9152# a_18_8152# w_n112_n8016#
+ a_n76_n500# w_n112_5580# w_n112_8052# a_18_n6680# a_n76_n2972# a_18_1972# a_n76_3208#
+ a_n76_n5444# a_18_4444# a_n76_6916# w_n112_n1836# a_18_n9152# a_n33_6819# w_n112_n4308#
+ VSUBS
X0 a_18_3208# a_n33_3111# a_n76_3208# w_n112_3108# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X1 a_18_n6680# a_n33_n6777# a_n76_n6680# w_n112_n6780# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X2 a_18_n500# a_n33_n597# a_n76_n500# w_n112_n600# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X3 a_18_n9152# a_n33_n9249# a_n76_n9152# w_n112_n9252# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X4 a_18_736# a_n33_639# a_n76_736# w_n112_636# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X5 a_18_n2972# a_n33_n3069# a_n76_n2972# w_n112_n3072# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X6 a_18_n7916# a_n33_n8013# a_n76_n7916# w_n112_n8016# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X7 a_18_5680# a_n33_5583# a_n76_5680# w_n112_5580# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X8 a_18_n5444# a_n33_n5541# a_n76_n5444# w_n112_n5544# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X9 a_18_8152# a_n33_8055# a_n76_8152# w_n112_8052# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X10 a_18_n1736# a_n33_n1833# a_n76_n1736# w_n112_n1836# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X11 a_18_6916# a_n33_6819# a_n76_6916# w_n112_6816# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X12 a_18_1972# a_n33_1875# a_n76_1972# w_n112_1872# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X13 a_18_n4208# a_n33_n4305# a_n76_n4208# w_n112_n4308# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X14 a_18_4444# a_n33_4347# a_n76_4444# w_n112_4344# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
C0 w_n112_8052# a_n33_8055# 0.106f
C1 a_n33_n597# a_18_n500# 0.0417f
C2 a_18_736# w_n112_n600# 0.00199f
C3 a_n33_n3069# w_n112_n1836# 4.13e-19
C4 a_18_n500# w_n112_636# 0.00199f
C5 a_n76_n5444# a_n33_n4305# 1.15e-19
C6 w_n112_n4308# a_n76_n2972# 0.00199f
C7 w_n112_n3072# a_18_n2972# 0.0182f
C8 a_n33_639# a_n76_n500# 1.15e-19
C9 a_n76_736# a_n33_n597# 1.15e-19
C10 a_n76_736# w_n112_636# 0.0182f
C11 a_n33_n1833# a_18_n1736# 0.0417f
C12 a_18_n1736# w_n112_n600# 0.00199f
C13 a_n33_n6777# w_n112_n6780# 0.106f
C14 a_n76_736# w_n112_1872# 0.00199f
C15 a_n76_n5444# a_n33_n6777# 1.15e-19
C16 a_n76_n500# w_n112_n1836# 0.00199f
C17 a_n76_n5444# w_n112_n4308# 0.00199f
C18 a_18_3208# a_n33_4347# 1.15e-19
C19 w_n112_n1836# a_18_n2972# 0.00199f
C20 a_n76_4444# a_18_4444# 0.747f
C21 a_n33_4347# a_n33_3111# 0.0665f
C22 w_n112_5580# a_n33_5583# 0.106f
C23 w_n112_6816# a_n33_8055# 4.13e-19
C24 a_n33_5583# a_18_5680# 0.0417f
C25 a_n33_n8013# a_18_n7916# 0.0417f
C26 w_n112_1872# a_n76_3208# 0.00199f
C27 w_n112_6816# a_n33_5583# 4.13e-19
C28 a_n33_639# a_n33_1875# 0.0665f
C29 w_n112_8052# a_n76_8152# 0.0182f
C30 a_n76_n500# a_18_n500# 0.747f
C31 a_n33_n597# a_n33_n1833# 0.0665f
C32 a_n33_n597# w_n112_n600# 0.106f
C33 w_n112_4344# a_n33_5583# 4.13e-19
C34 w_n112_n3072# a_n33_n4305# 4.13e-19
C35 a_18_n6680# w_n112_n6780# 0.0182f
C36 a_n76_n6680# w_n112_n8016# 0.00199f
C37 a_n76_3208# a_18_3208# 0.747f
C38 a_18_736# a_n33_n597# 1.15e-19
C39 a_n76_736# a_n76_n500# 0.00947f
C40 a_18_736# w_n112_636# 0.0182f
C41 a_18_n5444# w_n112_n5544# 0.0182f
C42 a_n76_3208# a_n33_3111# 0.0417f
C43 a_n33_n1833# a_n33_n3069# 0.0665f
C44 a_n33_n4305# a_n76_n4208# 0.0417f
C45 a_18_736# w_n112_1872# 0.00199f
C46 a_n76_4444# a_n33_3111# 1.15e-19
C47 w_n112_5580# a_n76_5680# 0.0182f
C48 a_n33_n597# a_18_n1736# 1.15e-19
C49 w_n112_6816# a_n76_8152# 0.00199f
C50 a_n33_5583# a_n33_4347# 0.0665f
C51 a_n76_5680# a_18_5680# 0.747f
C52 w_n112_n6780# a_n33_n5541# 4.13e-19
C53 a_n33_n8013# a_n33_n9249# 0.0665f
C54 w_n112_6816# a_n76_5680# 0.00199f
C55 a_n76_736# a_n33_1875# 1.15e-19
C56 a_n76_n5444# a_n33_n5541# 0.0417f
C57 a_n33_639# a_n76_1972# 1.15e-19
C58 w_n112_n4308# a_n76_n4208# 0.0182f
C59 w_n112_n3072# a_18_n4208# 0.00199f
C60 w_n112_n5544# a_n33_n4305# 4.13e-19
C61 w_n112_8052# a_18_8152# 0.0182f
C62 a_n76_n500# a_n33_n1833# 1.15e-19
C63 a_n76_n500# w_n112_n600# 0.0182f
C64 w_n112_4344# a_n76_5680# 0.00199f
C65 a_n76_n1736# a_n76_n2972# 0.00947f
C66 a_n33_n1833# a_18_n2972# 1.15e-19
C67 a_18_n1736# a_n33_n3069# 1.15e-19
C68 w_n112_3108# a_n33_4347# 4.13e-19
C69 a_n76_n4208# a_18_n4208# 0.747f
C70 a_n33_n8013# w_n112_n6780# 4.13e-19
C71 a_n76_3208# a_n33_1875# 1.15e-19
C72 a_n33_n6777# a_n76_n6680# 0.0417f
C73 a_n33_n597# w_n112_636# 4.13e-19
C74 a_n33_n6777# w_n112_n5544# 4.13e-19
C75 a_n33_n8013# a_18_n9152# 1.15e-19
C76 a_18_3208# a_18_4444# 0.00947f
C77 a_18_n7916# a_n33_n9249# 1.15e-19
C78 a_n76_n7916# a_n76_n9152# 0.00947f
C79 w_n112_n5544# a_18_n4208# 0.00199f
C80 a_18_4444# a_n33_3111# 1.15e-19
C81 w_n112_6816# a_18_8152# 0.00199f
C82 a_n33_5583# a_n76_4444# 1.15e-19
C83 a_n76_5680# a_n33_4347# 1.15e-19
C84 w_n112_3108# a_n76_3208# 0.0182f
C85 a_18_n1736# a_18_n2972# 0.00947f
C86 a_n76_736# a_n76_1972# 0.00947f
C87 a_n33_639# a_18_1972# 1.15e-19
C88 a_18_736# a_n33_1875# 1.15e-19
C89 a_n76_6916# a_18_6916# 0.747f
C90 w_n112_8052# a_n33_6819# 4.13e-19
C91 a_n33_n8013# w_n112_n9252# 4.13e-19
C92 a_n76_n6680# a_18_n6680# 0.747f
C93 w_n112_n6780# a_18_n7916# 0.00199f
C94 w_n112_n8016# a_n76_n7916# 0.0182f
C95 w_n112_1872# a_18_3208# 0.00199f
C96 a_18_n6680# w_n112_n5544# 0.00199f
C97 w_n112_3108# a_n76_4444# 0.00199f
C98 a_n76_n4208# a_n33_n5541# 1.15e-19
C99 w_n112_1872# a_n33_3111# 4.13e-19
C100 a_n76_3208# a_n76_1972# 0.00947f
C101 a_n33_n597# a_n76_n500# 0.0417f
C102 a_n76_n500# w_n112_636# 0.00199f
C103 a_18_n7916# a_18_n9152# 0.00947f
C104 a_n76_n1736# w_n112_n3072# 0.00199f
C105 a_18_3208# a_n33_3111# 0.0417f
C106 w_n112_5580# a_n33_6819# 4.13e-19
C107 a_n76_n6680# a_n33_n5541# 1.15e-19
C108 a_n33_6819# a_18_5680# 1.15e-19
C109 w_n112_n5544# a_n33_n5541# 0.106f
C110 w_n112_6816# a_n33_6819# 0.106f
C111 a_n76_6916# a_n33_8055# 1.15e-19
C112 a_n76_5680# a_n76_4444# 0.00947f
C113 a_n33_5583# a_18_4444# 1.15e-19
C114 a_n33_n3069# a_18_n2972# 0.0417f
C115 w_n112_n9252# a_18_n7916# 0.00199f
C116 a_n76_6916# a_n33_5583# 1.15e-19
C117 w_n112_636# a_n33_1875# 4.13e-19
C118 a_n76_n6680# a_n33_n8013# 1.15e-19
C119 a_n76_n1736# w_n112_n1836# 0.0182f
C120 w_n112_1872# a_n33_1875# 0.106f
C121 a_n33_n6777# a_n76_n7916# 1.15e-19
C122 w_n112_3108# a_18_4444# 0.00199f
C123 a_n33_n9249# a_18_n9152# 0.0417f
C124 a_18_3208# a_n33_1875# 1.15e-19
C125 a_n76_n5444# w_n112_n6780# 0.00199f
C126 a_n33_1875# a_n33_3111# 0.0665f
C127 a_18_6916# a_n33_8055# 1.15e-19
C128 a_n76_6916# a_n76_8152# 0.00947f
C129 w_n112_n8016# a_n76_n9152# 0.00199f
C130 w_n112_n9252# a_n33_n9249# 0.106f
C131 a_n33_n3069# a_n33_n4305# 0.0665f
C132 a_18_736# a_18_1972# 0.00947f
C133 a_n76_6916# a_n76_5680# 0.00947f
C134 a_18_6916# a_n33_5583# 1.15e-19
C135 w_n112_636# a_n76_1972# 0.00199f
C136 w_n112_3108# a_18_3208# 0.0182f
C137 w_n112_1872# a_n76_1972# 0.0182f
C138 w_n112_3108# a_n33_3111# 0.106f
C139 w_n112_n3072# a_n76_n2972# 0.0182f
C140 a_n33_n3069# w_n112_n4308# 4.13e-19
C141 a_n33_n1833# a_n76_n1736# 0.0417f
C142 a_n76_n1736# w_n112_n600# 0.00199f
C143 a_18_n2972# a_n33_n4305# 1.15e-19
C144 a_n76_n2972# a_n76_n4208# 0.00947f
C145 a_n76_1972# a_n33_3111# 1.15e-19
C146 w_n112_n9252# a_18_n9152# 0.0182f
C147 a_n33_n3069# a_18_n4208# 1.15e-19
C148 w_n112_n1836# a_n76_n2972# 0.00199f
C149 a_n33_n8013# a_n76_n7916# 0.0417f
C150 w_n112_636# a_18_1972# 0.00199f
C151 a_n76_n5444# a_n76_n4208# 0.00947f
C152 a_18_n5444# a_n33_n4305# 1.15e-19
C153 w_n112_n4308# a_18_n2972# 0.00199f
C154 w_n112_3108# a_n33_1875# 4.13e-19
C155 w_n112_1872# a_18_1972# 0.0182f
C156 a_n76_n1736# a_18_n1736# 0.747f
C157 a_18_n2972# a_18_n4208# 0.00947f
C158 a_n76_n6680# w_n112_n6780# 0.0182f
C159 a_n33_n6777# w_n112_n8016# 4.13e-19
C160 a_18_n5444# a_n33_n6777# 1.15e-19
C161 a_n76_n5444# a_n76_n6680# 0.00947f
C162 a_n76_n5444# w_n112_n5544# 0.0182f
C163 a_18_n5444# w_n112_n4308# 0.00199f
C164 a_n33_1875# a_n76_1972# 0.0417f
C165 a_18_3208# a_18_1972# 0.00947f
C166 w_n112_5580# a_18_5680# 0.0182f
C167 a_18_1972# a_n33_3111# 1.15e-19
C168 a_n33_8055# a_n76_8152# 0.0417f
C169 w_n112_6816# a_18_5680# 0.00199f
C170 a_18_n5444# a_18_n4208# 0.00947f
C171 a_n76_n7916# a_18_n7916# 0.747f
C172 a_n76_6916# a_n33_6819# 0.0417f
C173 a_18_6916# a_18_8152# 0.00947f
C174 a_n33_n597# a_n76_n1736# 1.15e-19
C175 w_n112_4344# a_18_5680# 0.00199f
C176 a_n33_5583# a_n76_5680# 0.0417f
C177 w_n112_n3072# a_n76_n4208# 0.00199f
C178 w_n112_n4308# a_n33_n4305# 0.106f
C179 w_n112_3108# a_n76_1972# 0.00199f
C180 a_18_n6680# w_n112_n8016# 0.00199f
C181 a_n33_n1833# a_n76_n2972# 1.15e-19
C182 a_18_n5444# a_18_n6680# 0.00947f
C183 a_n76_n1736# a_n33_n3069# 1.15e-19
C184 a_n33_n4305# a_18_n4208# 0.0417f
C185 a_n33_1875# a_18_1972# 0.0417f
C186 w_n112_5580# a_n33_4347# 4.13e-19
C187 a_18_5680# a_n33_4347# 1.15e-19
C188 a_n33_8055# a_18_8152# 0.0417f
C189 a_n33_n8013# a_n76_n9152# 1.15e-19
C190 a_18_n5444# a_n33_n5541# 0.0417f
C191 a_n76_n7916# a_n33_n9249# 1.15e-19
C192 w_n112_n5544# a_n76_n4208# 0.00199f
C193 w_n112_n4308# a_18_n4208# 0.0182f
C194 a_18_6916# a_n33_6819# 0.0417f
C195 a_n76_n500# a_n76_n1736# 0.00947f
C196 w_n112_4344# a_n33_4347# 0.106f
C197 a_n33_639# a_18_n500# 1.15e-19
C198 w_n112_3108# a_18_1972# 0.00199f
C199 a_n33_n8013# w_n112_n8016# 0.106f
C200 a_n33_n6777# a_18_n6680# 0.0417f
C201 w_n112_n6780# a_n76_n7916# 0.00199f
C202 a_18_n500# w_n112_n1836# 0.00199f
C203 a_n76_n6680# w_n112_n5544# 0.00199f
C204 a_n33_639# a_n76_736# 0.0417f
C205 a_n33_n4305# a_n33_n5541# 0.0665f
C206 w_n112_4344# a_n76_3208# 0.00199f
C207 a_n76_1972# a_18_1972# 0.747f
C208 w_n112_5580# a_n76_4444# 0.00199f
C209 a_n33_n1833# w_n112_n3072# 4.13e-19
C210 a_n76_8152# a_18_8152# 0.747f
C211 a_n33_8055# a_n33_6819# 0.0665f
C212 a_n33_n6777# a_n33_n5541# 0.0665f
C213 a_n33_5583# a_n33_6819# 0.0665f
C214 w_n112_n4308# a_n33_n5541# 4.13e-19
C215 w_n112_4344# a_n76_4444# 0.0182f
C216 a_n33_639# w_n112_n600# 4.13e-19
C217 w_n112_n8016# a_18_n7916# 0.0182f
C218 w_n112_n9252# a_n76_n7916# 0.00199f
C219 a_n33_n3069# a_n76_n2972# 0.0417f
C220 w_n112_8052# a_n76_6916# 0.00199f
C221 a_18_n4208# a_n33_n5541# 1.15e-19
C222 a_n33_n6777# a_n33_n8013# 0.0665f
C223 a_n33_n1833# w_n112_n1836# 0.106f
C224 a_n33_639# a_18_736# 0.0417f
C225 a_n76_3208# a_n33_4347# 1.15e-19
C226 a_18_n1736# w_n112_n3072# 0.00199f
C227 a_18_n6680# a_n33_n5541# 1.15e-19
C228 a_n33_n9249# a_n76_n9152# 0.0417f
C229 w_n112_5580# a_18_4444# 0.00199f
C230 a_18_n500# a_n33_n1833# 1.15e-19
C231 a_18_n500# w_n112_n600# 0.0182f
C232 a_n76_n2972# a_18_n2972# 0.747f
C233 a_n33_4347# a_n76_4444# 0.0417f
C234 a_18_5680# a_18_4444# 0.00947f
C235 w_n112_5580# a_n76_6916# 0.00199f
C236 a_n76_8152# a_n33_6819# 1.15e-19
C237 a_n76_5680# a_n33_6819# 1.15e-19
C238 w_n112_4344# a_18_4444# 0.0182f
C239 w_n112_6816# a_n76_6916# 0.0182f
C240 a_18_736# a_18_n500# 0.00947f
C241 a_n76_736# w_n112_n600# 0.00199f
C242 a_18_n6680# a_n33_n8013# 1.15e-19
C243 w_n112_n8016# a_n33_n9249# 4.13e-19
C244 a_18_n1736# w_n112_n1836# 0.0182f
C245 a_n76_n6680# a_n76_n7916# 0.00947f
C246 a_n33_n6777# a_18_n7916# 1.15e-19
C247 w_n112_8052# a_18_6916# 0.00199f
C248 a_n33_639# a_n33_n597# 0.0665f
C249 a_n76_736# a_18_736# 0.747f
C250 a_n33_639# w_n112_636# 0.106f
C251 a_n76_n9152# a_18_n9152# 0.747f
C252 a_n76_3208# a_n76_4444# 0.00947f
C253 a_18_n500# a_18_n1736# 0.00947f
C254 a_18_n5444# w_n112_n6780# 0.00199f
C255 a_n33_n3069# w_n112_n3072# 0.106f
C256 a_n33_639# w_n112_1872# 4.13e-19
C257 a_n76_n5444# a_18_n5444# 0.747f
C258 a_n33_n597# w_n112_n1836# 4.13e-19
C259 a_n33_n1833# w_n112_n600# 4.13e-19
C260 a_n76_n2972# a_n33_n4305# 1.15e-19
C261 a_n33_4347# a_18_4444# 0.0417f
C262 w_n112_5580# a_18_6916# 0.00199f
C263 a_18_8152# a_n33_6819# 1.15e-19
C264 w_n112_4344# a_18_3208# 0.00199f
C265 w_n112_n9252# a_n76_n9152# 0.0182f
C266 w_n112_n8016# a_18_n9152# 0.00199f
C267 a_n33_n3069# a_n76_n4208# 1.15e-19
C268 a_18_6916# a_18_5680# 0.00947f
C269 a_18_n6680# a_18_n7916# 0.00947f
C270 w_n112_4344# a_n33_3111# 4.13e-19
C271 w_n112_6816# a_18_6916# 0.0182f
C272 a_18_n9152# VSUBS 0.426f
C273 a_n76_n9152# VSUBS 0.426f
C274 a_n33_n9249# VSUBS 0.192f
C275 a_18_n7916# VSUBS 0.415f
C276 a_n76_n7916# VSUBS 0.415f
C277 a_n33_n8013# VSUBS 0.156f
C278 a_18_n6680# VSUBS 0.415f
C279 a_n76_n6680# VSUBS 0.415f
C280 a_n33_n6777# VSUBS 0.156f
C281 a_18_n5444# VSUBS 0.415f
C282 a_n76_n5444# VSUBS 0.415f
C283 a_n33_n5541# VSUBS 0.156f
C284 a_18_n4208# VSUBS 0.415f
C285 a_n76_n4208# VSUBS 0.415f
C286 a_n33_n4305# VSUBS 0.156f
C287 a_18_n2972# VSUBS 0.415f
C288 a_n76_n2972# VSUBS 0.415f
C289 a_n33_n3069# VSUBS 0.156f
C290 a_18_n1736# VSUBS 0.415f
C291 a_n76_n1736# VSUBS 0.415f
C292 a_n33_n1833# VSUBS 0.156f
C293 a_18_n500# VSUBS 0.415f
C294 a_n76_n500# VSUBS 0.415f
C295 a_n33_n597# VSUBS 0.156f
C296 a_18_736# VSUBS 0.415f
C297 a_n76_736# VSUBS 0.415f
C298 a_n33_639# VSUBS 0.156f
C299 a_18_1972# VSUBS 0.415f
C300 a_n76_1972# VSUBS 0.415f
C301 a_n33_1875# VSUBS 0.156f
C302 a_18_3208# VSUBS 0.415f
C303 a_n76_3208# VSUBS 0.415f
C304 a_n33_3111# VSUBS 0.156f
C305 a_18_4444# VSUBS 0.415f
C306 a_n76_4444# VSUBS 0.415f
C307 a_n33_4347# VSUBS 0.156f
C308 a_18_5680# VSUBS 0.415f
C309 a_n76_5680# VSUBS 0.415f
C310 a_n33_5583# VSUBS 0.156f
C311 a_18_6916# VSUBS 0.415f
C312 a_n76_6916# VSUBS 0.415f
C313 a_n33_6819# VSUBS 0.156f
C314 a_18_8152# VSUBS 0.426f
C315 a_n76_8152# VSUBS 0.426f
C316 a_n33_8055# VSUBS 0.192f
C317 w_n112_n9252# VSUBS 0.806f
C318 w_n112_n8016# VSUBS 0.806f
C319 w_n112_n6780# VSUBS 0.806f
C320 w_n112_n5544# VSUBS 0.806f
C321 w_n112_n4308# VSUBS 0.806f
C322 w_n112_n3072# VSUBS 0.806f
C323 w_n112_n1836# VSUBS 0.806f
C324 w_n112_n600# VSUBS 0.806f
C325 w_n112_636# VSUBS 0.806f
C326 w_n112_1872# VSUBS 0.806f
C327 w_n112_3108# VSUBS 0.806f
C328 w_n112_4344# VSUBS 0.806f
C329 w_n112_5580# VSUBS 0.806f
C330 w_n112_6816# VSUBS 0.806f
C331 w_n112_8052# VSUBS 0.806f
.ends

.subckt sky130_fd_pr__nfet_01v8_MHE452 a_n158_n359# a_n100_957# a_100_n1295# a_n158_577#
+ a_n100_21# a_100_109# a_n100_n915# a_100_n827# a_n100_489# a_100_1045# a_n158_n1295#
+ a_n158_n827# a_100_577# a_n158_1045# a_n100_n447# a_n158_109# a_100_n359# a_n100_n1383#
+ VSUBS
X0 a_100_n827# a_n100_n915# a_n158_n827# VSUBS sky130_fd_pr__nfet_01v8 ad=0.363 pd=3.08 as=0.363 ps=3.08 w=1.25 l=1
**devattr s=14500,616 d=14500,616
X1 a_100_n359# a_n100_n447# a_n158_n359# VSUBS sky130_fd_pr__nfet_01v8 ad=0.363 pd=3.08 as=0.363 ps=3.08 w=1.25 l=1
**devattr s=14500,616 d=14500,616
X2 a_100_577# a_n100_489# a_n158_577# VSUBS sky130_fd_pr__nfet_01v8 ad=0.363 pd=3.08 as=0.363 ps=3.08 w=1.25 l=1
**devattr s=14500,616 d=14500,616
X3 a_100_1045# a_n100_957# a_n158_1045# VSUBS sky130_fd_pr__nfet_01v8 ad=0.363 pd=3.08 as=0.363 ps=3.08 w=1.25 l=1
**devattr s=14500,616 d=14500,616
X4 a_100_n1295# a_n100_n1383# a_n158_n1295# VSUBS sky130_fd_pr__nfet_01v8 ad=0.363 pd=3.08 as=0.363 ps=3.08 w=1.25 l=1
**devattr s=14500,616 d=14500,616
X5 a_100_109# a_n100_21# a_n158_109# VSUBS sky130_fd_pr__nfet_01v8 ad=0.363 pd=3.08 as=0.363 ps=3.08 w=1.25 l=1
**devattr s=14500,616 d=14500,616
C0 a_n158_109# a_n158_577# 0.0113f
C1 a_100_n827# a_100_n359# 0.0113f
C2 a_n100_n447# a_n158_n359# 0.0322f
C3 a_n100_957# a_100_1045# 0.0322f
C4 a_n100_n915# a_n100_n1383# 0.205f
C5 a_100_n359# a_n100_n447# 0.0322f
C6 a_100_n827# a_n100_n915# 0.0322f
C7 a_n100_n915# a_n100_n447# 0.205f
C8 a_n100_957# a_n100_489# 0.205f
C9 a_n158_1045# a_n158_577# 0.0113f
C10 a_n158_n1295# a_n100_n1383# 0.0322f
C11 a_100_1045# a_100_577# 0.0113f
C12 a_n100_21# a_n100_489# 0.205f
C13 a_n100_489# a_100_577# 0.0322f
C14 a_n100_21# a_100_109# 0.0322f
C15 a_100_109# a_100_577# 0.0113f
C16 a_n158_n359# a_n158_n827# 0.0113f
C17 a_100_109# a_n158_109# 0.0693f
C18 a_n100_21# a_n158_109# 0.0322f
C19 a_100_n359# a_100_109# 0.0113f
C20 a_n100_957# a_n158_1045# 0.0322f
C21 a_n100_n915# a_n158_n827# 0.0322f
C22 a_n158_109# a_n158_n359# 0.0113f
C23 a_n158_1045# a_100_1045# 0.0693f
C24 a_100_n359# a_n158_n359# 0.0693f
C25 a_n158_n1295# a_n158_n827# 0.0113f
C26 a_n158_n1295# a_100_n1295# 0.0693f
C27 a_n100_489# a_n158_577# 0.0322f
C28 a_100_n827# a_n158_n827# 0.0693f
C29 a_100_n1295# a_n100_n1383# 0.0322f
C30 a_n158_577# a_100_577# 0.0693f
C31 a_100_n827# a_100_n1295# 0.0113f
C32 a_n100_21# a_n100_n447# 0.205f
C33 a_100_n1295# VSUBS 0.14f
C34 a_n158_n1295# VSUBS 0.14f
C35 a_n100_n1383# VSUBS 0.553f
C36 a_100_n827# VSUBS 0.13f
C37 a_n158_n827# VSUBS 0.13f
C38 a_n100_n915# VSUBS 0.441f
C39 a_100_n359# VSUBS 0.13f
C40 a_n158_n359# VSUBS 0.13f
C41 a_n100_n447# VSUBS 0.441f
C42 a_100_109# VSUBS 0.13f
C43 a_n158_109# VSUBS 0.13f
C44 a_n100_21# VSUBS 0.441f
C45 a_100_577# VSUBS 0.13f
C46 a_n158_577# VSUBS 0.13f
C47 a_n100_489# VSUBS 0.441f
C48 a_100_1045# VSUBS 0.14f
C49 a_n158_1045# VSUBS 0.14f
C50 a_n100_957# VSUBS 0.553f
.ends

.subckt sky130_fd_pr__pfet_01v8_P2UXFR a_n300_n1215# w_n394_n1218# a_n358_n1118# a_n300_21#
+ a_300_118# w_n394_18# a_300_n1118# a_n358_118# VSUBS
X0 a_300_118# a_n300_21# a_n358_118# w_n394_18# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=3
**devattr s=58000,2116 d=58000,2116
X1 a_300_n1118# a_n300_n1215# a_n358_n1118# w_n394_n1218# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=3
**devattr s=58000,2116 d=58000,2116
C0 a_n358_118# a_n358_n1118# 0.0105f
C1 w_n394_18# a_n358_118# 0.0187f
C2 a_n300_21# w_n394_18# 0.382f
C3 a_300_118# a_300_n1118# 0.0105f
C4 a_300_118# a_n358_118# 0.107f
C5 a_n300_21# a_300_118# 0.184f
C6 a_n300_n1215# w_n394_n1218# 0.382f
C7 a_n300_21# a_n358_118# 0.184f
C8 a_n358_n1118# w_n394_n1218# 0.0187f
C9 a_n300_n1215# a_n358_n1118# 0.184f
C10 w_n394_18# a_n300_n1215# 0.00346f
C11 w_n394_18# a_n358_n1118# 0.0023f
C12 a_300_n1118# w_n394_n1218# 0.0187f
C13 a_300_118# w_n394_n1218# 0.0023f
C14 a_n300_n1215# a_300_n1118# 0.184f
C15 a_300_n1118# a_n358_n1118# 0.107f
C16 a_n358_118# w_n394_n1218# 0.0023f
C17 a_n300_21# w_n394_n1218# 0.00346f
C18 w_n394_18# a_300_n1118# 0.0023f
C19 a_n300_21# a_n300_n1215# 0.62f
C20 w_n394_18# a_300_118# 0.0187f
C21 a_300_n1118# VSUBS 0.536f
C22 a_n358_n1118# VSUBS 0.536f
C23 a_n300_n1215# VSUBS 1.08f
C24 a_300_118# VSUBS 0.536f
C25 a_n358_118# VSUBS 0.536f
C26 a_n300_21# VSUBS 1.08f
C27 w_n394_n1218# VSUBS 2.84f
C28 w_n394_18# VSUBS 2.84f
.ends

.subckt sky130_fd_pr__pfet_01v8_MGA63L a_18_n500# a_n33_n597# w_n112_n600# a_n76_n500#
+ VSUBS
X0 a_18_n500# a_n33_n597# a_n76_n500# w_n112_n600# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
C0 a_n76_n500# w_n112_n600# 0.0182f
C1 a_n76_n500# a_18_n500# 0.747f
C2 a_18_n500# w_n112_n600# 0.0182f
C3 a_n76_n500# a_n33_n597# 0.0417f
C4 a_n33_n597# w_n112_n600# 0.106f
C5 a_18_n500# a_n33_n597# 0.0417f
C6 a_18_n500# VSUBS 0.437f
C7 a_n76_n500# VSUBS 0.437f
C8 a_n33_n597# VSUBS 0.228f
C9 w_n112_n600# VSUBS 0.806f
.ends

.subckt sky130_fd_pr__nfet_01v8_VT3ZQW a_n158_n125# a_n100_n213# a_100_n125# VSUBS
X0 a_100_n125# a_n100_n213# a_n158_n125# VSUBS sky130_fd_pr__nfet_01v8 ad=0.363 pd=3.08 as=0.363 ps=3.08 w=1.25 l=1
**devattr s=14500,616 d=14500,616
C0 a_100_n125# a_n100_n213# 0.0322f
C1 a_100_n125# a_n158_n125# 0.0693f
C2 a_n158_n125# a_n100_n213# 0.0322f
C3 a_100_n125# VSUBS 0.151f
C4 a_n158_n125# VSUBS 0.151f
C5 a_n100_n213# VSUBS 0.664f
.ends

.subckt sky130_fd_pr__pfet_01v8_RRUZAE a_n358_n2972# a_n300_n1833# a_n300_n3069# w_n394_n1836#
+ w_n394_1872# a_n358_n1736# a_300_736# a_300_1972# a_300_n2972# w_n394_636# w_n394_n3072#
+ a_n300_n597# a_300_n500# a_n300_639# a_n358_1972# a_n300_1875# w_n394_n600# a_300_n1736#
+ a_n358_n500# a_n358_736# VSUBS
X0 a_300_n500# a_n300_n597# a_n358_n500# w_n394_n600# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=3
**devattr s=58000,2116 d=58000,2116
X1 a_300_736# a_n300_639# a_n358_736# w_n394_636# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=3
**devattr s=58000,2116 d=58000,2116
X2 a_300_n2972# a_n300_n3069# a_n358_n2972# w_n394_n3072# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=3
**devattr s=58000,2116 d=58000,2116
X3 a_300_1972# a_n300_1875# a_n358_1972# w_n394_1872# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=3
**devattr s=58000,2116 d=58000,2116
X4 a_300_n1736# a_n300_n1833# a_n358_n1736# w_n394_n1836# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=3
**devattr s=58000,2116 d=58000,2116
C0 a_n358_1972# w_n394_1872# 0.0187f
C1 a_300_n2972# a_n300_n3069# 0.184f
C2 a_300_1972# a_n358_1972# 0.107f
C3 a_300_736# w_n394_1872# 0.0023f
C4 w_n394_n600# a_n358_n500# 0.0187f
C5 w_n394_n1836# a_n300_n3069# 0.00346f
C6 a_300_736# a_300_1972# 0.0105f
C7 a_n300_1875# w_n394_1872# 0.382f
C8 a_n358_n1736# a_300_n1736# 0.107f
C9 a_300_1972# a_n300_1875# 0.184f
C10 a_300_736# a_n300_639# 0.184f
C11 w_n394_n1836# a_n358_n500# 0.0023f
C12 a_300_n500# w_n394_636# 0.0023f
C13 a_300_n500# a_300_n1736# 0.0105f
C14 a_n358_n1736# a_n358_n2972# 0.0105f
C15 a_n300_639# a_n300_1875# 0.62f
C16 a_n358_n1736# a_n300_n1833# 0.184f
C17 a_300_n1736# a_n300_n1833# 0.184f
C18 a_n358_1972# w_n394_636# 0.0023f
C19 a_300_736# w_n394_636# 0.0187f
C20 a_n300_1875# w_n394_636# 0.00346f
C21 a_300_736# a_300_n500# 0.0105f
C22 w_n394_n600# a_n300_n597# 0.382f
C23 a_n358_n1736# a_n358_n500# 0.0105f
C24 w_n394_636# a_n358_n500# 0.0023f
C25 a_n358_n2972# a_n300_n3069# 0.184f
C26 w_n394_n600# a_n358_736# 0.0023f
C27 a_n300_n1833# a_n300_n3069# 0.62f
C28 a_300_n500# a_n358_n500# 0.107f
C29 a_n300_n597# w_n394_n1836# 0.00346f
C30 a_n358_1972# a_n300_1875# 0.184f
C31 w_n394_n3072# a_300_n2972# 0.0187f
C32 w_n394_1872# a_n358_736# 0.0023f
C33 a_n300_n597# a_n300_639# 0.62f
C34 a_n300_639# a_n358_736# 0.184f
C35 w_n394_n1836# a_300_n2972# 0.0023f
C36 w_n394_n600# a_n300_639# 0.00346f
C37 a_300_1972# w_n394_1872# 0.0187f
C38 a_n300_n597# w_n394_636# 0.00346f
C39 a_n300_639# w_n394_1872# 0.00346f
C40 a_n300_n597# a_300_n500# 0.184f
C41 w_n394_636# a_n358_736# 0.0187f
C42 a_n358_n1736# w_n394_n3072# 0.0023f
C43 w_n394_n600# a_n358_n1736# 0.0023f
C44 w_n394_n3072# a_300_n1736# 0.0023f
C45 a_n300_n597# a_n300_n1833# 0.62f
C46 w_n394_n600# a_300_n1736# 0.0023f
C47 w_n394_n600# a_300_n500# 0.0187f
C48 a_300_n1736# a_300_n2972# 0.0105f
C49 a_n358_n2972# w_n394_n3072# 0.0187f
C50 a_n358_n1736# w_n394_n1836# 0.0187f
C51 w_n394_n3072# a_n300_n1833# 0.00346f
C52 a_300_n1736# w_n394_n1836# 0.0187f
C53 w_n394_n600# a_n300_n1833# 0.00346f
C54 a_n358_1972# a_n358_736# 0.0105f
C55 a_300_1972# w_n394_636# 0.0023f
C56 a_n358_n2972# a_300_n2972# 0.107f
C57 a_300_736# a_n358_736# 0.107f
C58 a_300_n500# w_n394_n1836# 0.0023f
C59 a_n358_n2972# w_n394_n1836# 0.0023f
C60 a_n300_n597# a_n358_n500# 0.184f
C61 a_n300_639# w_n394_636# 0.382f
C62 w_n394_n600# a_300_736# 0.0023f
C63 w_n394_n3072# a_n300_n3069# 0.382f
C64 w_n394_n1836# a_n300_n1833# 0.382f
C65 a_n358_n500# a_n358_736# 0.0105f
C66 a_300_n2972# VSUBS 0.536f
C67 a_n358_n2972# VSUBS 0.536f
C68 a_n300_n3069# VSUBS 1.08f
C69 a_300_n1736# VSUBS 0.524f
C70 a_n358_n1736# VSUBS 0.524f
C71 a_n300_n1833# VSUBS 0.739f
C72 a_300_n500# VSUBS 0.524f
C73 a_n358_n500# VSUBS 0.524f
C74 a_n300_n597# VSUBS 0.739f
C75 a_300_736# VSUBS 0.524f
C76 a_n358_736# VSUBS 0.524f
C77 a_n300_639# VSUBS 0.739f
C78 a_300_1972# VSUBS 0.536f
C79 a_n358_1972# VSUBS 0.536f
C80 a_n300_1875# VSUBS 1.08f
C81 w_n394_n3072# VSUBS 2.84f
C82 w_n394_n1836# VSUBS 2.84f
C83 w_n394_n600# VSUBS 2.84f
C84 w_n394_636# VSUBS 2.84f
C85 w_n394_1872# VSUBS 2.84f
.ends

.subckt sky130_fd_pr__pfet_01v8_8DHNHY w_n112_636# a_n33_n5541# a_n33_n8013# a_n76_736#
+ a_n33_9291# w_n112_1872# a_18_9388# w_n112_4344# a_18_n500# a_18_n2972# a_18_n5444#
+ a_n76_n1736# a_n33_3111# a_n76_n4208# a_18_3208# w_n112_9288# a_n76_n7916# a_n33_n1833#
+ a_18_6916# a_n76_5680# w_n112_n3072# a_n76_n10388# a_n33_n4305# a_n33_5583# a_n76_8152#
+ w_n112_n6780# a_n33_8055# a_n33_n3069# a_n33_639# w_n112_n9252# w_n112_3108# a_18_n10388#
+ w_n112_6816# a_n33_n6777# a_n33_n597# w_n112_n10488# a_n33_n9249# a_18_n1736# a_18_n4208#
+ a_18_n7916# a_n76_1972# a_n33_1875# w_n112_n600# a_n76_n6680# a_18_736# a_n76_4444#
+ a_18_5680# a_n33_4347# w_n112_n5544# a_n76_n9152# a_18_8152# w_n112_n8016# a_n76_n500#
+ a_n76_9388# w_n112_5580# w_n112_8052# a_18_n6680# a_n76_n2972# a_18_1972# a_n76_3208#
+ a_n76_n5444# a_18_4444# a_n76_6916# w_n112_n1836# a_n33_n10485# a_18_n9152# a_n33_6819#
+ w_n112_n4308# VSUBS
X0 a_18_3208# a_n33_3111# a_n76_3208# w_n112_3108# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X1 a_18_n6680# a_n33_n6777# a_n76_n6680# w_n112_n6780# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X2 a_18_9388# a_n33_9291# a_n76_9388# w_n112_9288# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X3 a_18_n500# a_n33_n597# a_n76_n500# w_n112_n600# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X4 a_18_n9152# a_n33_n9249# a_n76_n9152# w_n112_n9252# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X5 a_18_736# a_n33_639# a_n76_736# w_n112_636# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X6 a_18_n2972# a_n33_n3069# a_n76_n2972# w_n112_n3072# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X7 a_18_n7916# a_n33_n8013# a_n76_n7916# w_n112_n8016# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X8 a_18_5680# a_n33_5583# a_n76_5680# w_n112_5580# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X9 a_18_n5444# a_n33_n5541# a_n76_n5444# w_n112_n5544# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X10 a_18_8152# a_n33_8055# a_n76_8152# w_n112_8052# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X11 a_18_n1736# a_n33_n1833# a_n76_n1736# w_n112_n1836# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X12 a_18_6916# a_n33_6819# a_n76_6916# w_n112_6816# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X13 a_18_1972# a_n33_1875# a_n76_1972# w_n112_1872# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X14 a_18_n4208# a_n33_n4305# a_n76_n4208# w_n112_n4308# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X15 a_18_4444# a_n33_4347# a_n76_4444# w_n112_4344# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X16 a_18_n10388# a_n33_n10485# a_n76_n10388# w_n112_n10488# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
C0 w_n112_n5544# a_n33_n4305# 4.13e-19
C1 a_18_736# a_n33_1875# 1.15e-19
C2 a_18_736# w_n112_n600# 0.00199f
C3 w_n112_n4308# a_18_n4208# 0.0182f
C4 a_n33_6819# w_n112_5580# 4.13e-19
C5 a_18_n5444# w_n112_n6780# 0.00199f
C6 a_n76_736# w_n112_636# 0.0182f
C7 a_18_n10388# w_n112_n10488# 0.0182f
C8 a_18_1972# a_n33_1875# 0.0417f
C9 a_18_n6680# w_n112_n6780# 0.0182f
C10 w_n112_6816# a_n33_5583# 4.13e-19
C11 a_n76_n1736# a_n76_n2972# 0.00947f
C12 w_n112_4344# a_18_4444# 0.0182f
C13 a_n33_n1833# a_18_n2972# 1.15e-19
C14 a_18_n1736# a_n33_n3069# 1.15e-19
C15 a_n76_n500# a_18_n500# 0.747f
C16 a_18_5680# a_n76_5680# 0.747f
C17 w_n112_n5544# a_18_n4208# 0.00199f
C18 a_n33_n5541# a_n76_n5444# 0.0417f
C19 w_n112_8052# a_n33_9291# 4.13e-19
C20 a_18_4444# a_n33_3111# 1.15e-19
C21 w_n112_4344# a_n76_3208# 0.00199f
C22 a_n33_n8013# a_n33_n9249# 0.0665f
C23 a_18_5680# w_n112_5580# 0.0182f
C24 w_n112_n8016# a_18_n6680# 0.00199f
C25 a_n76_1972# a_n76_3208# 0.00947f
C26 a_n33_6819# a_n33_8055# 0.0665f
C27 a_n33_n597# w_n112_n600# 0.106f
C28 w_n112_n4308# a_n33_n5541# 4.13e-19
C29 w_n112_4344# a_n33_4347# 0.106f
C30 a_18_1972# w_n112_3108# 0.00199f
C31 a_n76_n6680# a_n33_n5541# 1.15e-19
C32 a_n33_3111# a_n76_3208# 0.0417f
C33 a_n33_n6777# w_n112_n6780# 0.106f
C34 w_n112_n3072# a_n33_n1833# 4.13e-19
C35 a_18_736# w_n112_636# 0.0182f
C36 w_n112_8052# a_n76_8152# 0.0182f
C37 w_n112_4344# a_n33_5583# 4.13e-19
C38 a_18_6916# a_n33_5583# 1.15e-19
C39 a_18_n1736# a_18_n2972# 0.00947f
C40 a_n33_4347# a_n33_3111# 0.0665f
C41 a_n33_9291# a_n76_8152# 1.15e-19
C42 a_n33_639# a_n33_1875# 0.0665f
C43 w_n112_n600# a_n33_639# 4.13e-19
C44 a_n33_n8013# w_n112_n6780# 4.13e-19
C45 w_n112_6816# a_n76_8152# 0.00199f
C46 a_18_1972# w_n112_636# 0.00199f
C47 a_n76_n5444# a_18_n5444# 0.747f
C48 w_n112_n8016# a_n33_n6777# 4.13e-19
C49 a_18_n7916# a_n33_n9249# 1.15e-19
C50 a_n76_n7916# a_n76_n9152# 0.00947f
C51 w_n112_n600# a_n76_n1736# 0.00199f
C52 w_n112_8052# a_18_6916# 0.00199f
C53 w_n112_8052# a_n76_9388# 0.00199f
C54 w_n112_n5544# a_n33_n5541# 0.106f
C55 w_n112_n1836# a_n33_n1833# 0.106f
C56 w_n112_n4308# a_18_n5444# 0.00199f
C57 a_n76_9388# a_n33_9291# 0.0417f
C58 a_18_4444# w_n112_5580# 0.00199f
C59 w_n112_n8016# a_n33_n8013# 0.106f
C60 a_18_9388# a_18_8152# 0.00947f
C61 w_n112_n3072# a_18_n1736# 0.00199f
C62 a_n33_n4305# a_n33_n3069# 0.0665f
C63 w_n112_6816# a_18_6916# 0.0182f
C64 w_n112_1872# a_n76_3208# 0.00199f
C65 a_n76_n500# w_n112_n600# 0.0182f
C66 a_n33_9291# w_n112_9288# 0.106f
C67 a_n33_n8013# w_n112_n9252# 4.13e-19
C68 a_n33_n597# w_n112_636# 4.13e-19
C69 a_n76_n6680# a_18_n6680# 0.747f
C70 a_18_n7916# w_n112_n6780# 0.00199f
C71 a_n33_4347# a_n76_5680# 1.15e-19
C72 a_18_n9152# a_n33_n10485# 1.15e-19
C73 a_n76_6916# a_n33_5583# 1.15e-19
C74 a_n33_n3069# a_18_n2972# 0.0417f
C75 a_n76_9388# a_n76_8152# 0.00947f
C76 a_n76_n9152# a_18_n9152# 0.747f
C77 a_n76_5680# a_n33_5583# 0.0417f
C78 a_n33_4347# w_n112_5580# 4.13e-19
C79 a_n33_639# w_n112_636# 0.106f
C80 w_n112_n5544# a_18_n5444# 0.0182f
C81 a_n76_n5444# a_n33_n6777# 1.15e-19
C82 a_n76_8152# w_n112_9288# 0.00199f
C83 a_n33_5583# w_n112_5580# 0.106f
C84 w_n112_n1836# a_18_n1736# 0.0182f
C85 w_n112_n8016# a_18_n7916# 0.0182f
C86 a_n33_n4305# a_18_n2972# 1.15e-19
C87 w_n112_8052# a_n76_6916# 0.00199f
C88 a_n76_n4208# a_n76_n2972# 0.00947f
C89 a_18_n4208# a_n33_n3069# 1.15e-19
C90 a_18_n6680# w_n112_n5544# 0.00199f
C91 a_n76_n6680# a_n33_n6777# 0.0417f
C92 w_n112_4344# a_n33_3111# 4.13e-19
C93 w_n112_n3072# a_n33_n3069# 0.106f
C94 a_18_n7916# w_n112_n9252# 0.00199f
C95 w_n112_6816# a_n76_6916# 0.0182f
C96 a_n76_1972# a_n33_3111# 1.15e-19
C97 a_18_n9152# a_18_n10388# 0.00947f
C98 w_n112_6816# a_n76_5680# 0.00199f
C99 a_18_n500# w_n112_n600# 0.0182f
C100 a_n76_9388# w_n112_9288# 0.0182f
C101 a_n33_n4305# a_18_n4208# 0.0417f
C102 a_n76_n500# w_n112_636# 0.00199f
C103 a_n76_n6680# a_n33_n8013# 1.15e-19
C104 a_n33_n597# a_n33_n1833# 0.0665f
C105 a_n76_6916# a_n76_8152# 0.00947f
C106 a_n33_n9249# a_n76_n10388# 1.15e-19
C107 a_n76_n9152# a_n33_n10485# 1.15e-19
C108 a_n33_n4305# w_n112_n3072# 4.13e-19
C109 a_18_3208# a_n33_1875# 1.15e-19
C110 a_18_n4208# a_18_n2972# 0.00947f
C111 w_n112_n5544# a_n33_n6777# 4.13e-19
C112 a_n33_6819# a_18_8152# 1.15e-19
C113 w_n112_n1836# a_n33_n3069# 4.13e-19
C114 a_n76_736# a_n76_1972# 0.00947f
C115 w_n112_n8016# a_n33_n9249# 4.13e-19
C116 w_n112_n3072# a_18_n2972# 0.0182f
C117 a_18_6916# a_n76_6916# 0.747f
C118 w_n112_4344# a_n76_5680# 0.00199f
C119 w_n112_8052# a_n33_8055# 0.106f
C120 w_n112_1872# a_n76_1972# 0.0182f
C121 a_n33_n1833# a_n76_n1736# 0.0417f
C122 a_n33_n9249# w_n112_n9252# 0.106f
C123 a_n33_9291# a_n33_8055# 0.0665f
C124 a_n33_n10485# a_18_n10388# 0.0417f
C125 a_n33_n597# a_18_n1736# 1.15e-19
C126 w_n112_1872# a_n33_3111# 4.13e-19
C127 w_n112_6816# a_n33_8055# 4.13e-19
C128 a_18_6916# w_n112_5580# 0.00199f
C129 a_18_n4208# w_n112_n3072# 0.00199f
C130 a_n33_n4305# a_n33_n5541# 0.0665f
C131 a_18_n500# w_n112_636# 0.00199f
C132 a_18_3208# w_n112_3108# 0.0182f
C133 a_n76_n500# a_n33_n1833# 1.15e-19
C134 a_n33_8055# a_n76_8152# 0.0417f
C135 w_n112_n1836# a_18_n2972# 0.00199f
C136 a_n76_n10388# w_n112_n9252# 0.00199f
C137 a_n76_n1736# a_18_n1736# 0.747f
C138 a_n76_n7916# a_n33_n6777# 1.15e-19
C139 a_n33_n9249# w_n112_n10488# 4.13e-19
C140 a_n76_4444# w_n112_3108# 0.00199f
C141 a_n76_736# w_n112_1872# 0.00199f
C142 w_n112_n4308# a_n76_n2972# 0.00199f
C143 a_n76_6916# a_n76_5680# 0.00947f
C144 a_18_6916# a_n33_8055# 1.15e-19
C145 a_n76_9388# a_n33_8055# 1.15e-19
C146 a_18_n4208# a_n33_n5541# 1.15e-19
C147 a_n76_n4208# a_n76_n5444# 0.00947f
C148 a_n33_n4305# a_18_n5444# 1.15e-19
C149 a_n33_n8013# a_n76_n7916# 0.0417f
C150 a_n76_1972# a_18_1972# 0.747f
C151 a_n76_6916# w_n112_5580# 0.00199f
C152 a_n76_5680# w_n112_5580# 0.0182f
C153 a_n33_8055# w_n112_9288# 4.13e-19
C154 w_n112_n4308# a_n76_n4208# 0.0182f
C155 a_n33_1875# w_n112_3108# 4.13e-19
C156 a_18_1972# a_n33_3111# 1.15e-19
C157 a_n76_n5444# w_n112_n6780# 0.00199f
C158 a_18_n500# a_n33_n1833# 1.15e-19
C159 a_n76_n10388# w_n112_n10488# 0.0182f
C160 a_n76_736# a_18_736# 0.747f
C161 a_n76_n6680# w_n112_n6780# 0.0182f
C162 a_n76_n1736# a_n33_n3069# 1.15e-19
C163 w_n112_636# a_n33_1875# 4.13e-19
C164 a_n33_n1833# a_n76_n2972# 1.15e-19
C165 a_n33_n8013# a_18_n9152# 1.15e-19
C166 a_18_n4208# a_18_n5444# 0.00947f
C167 a_18_736# w_n112_1872# 0.00199f
C168 a_n76_n7916# a_18_n7916# 0.747f
C169 a_n76_6916# a_n33_8055# 1.15e-19
C170 w_n112_n5544# a_n76_n4208# 0.00199f
C171 a_18_4444# a_18_3208# 0.00947f
C172 w_n112_n8016# a_n76_n6680# 0.00199f
C173 a_n76_1972# a_n33_639# 1.15e-19
C174 a_18_n500# a_18_n1736# 0.00947f
C175 w_n112_1872# a_18_1972# 0.0182f
C176 a_n76_3208# a_18_3208# 0.747f
C177 a_n76_4444# a_18_4444# 0.747f
C178 a_18_n7916# a_18_n9152# 0.00947f
C179 w_n112_8052# a_18_8152# 0.0182f
C180 a_n33_4347# a_18_3208# 1.15e-19
C181 a_n76_736# a_n33_n597# 1.15e-19
C182 a_18_8152# a_n33_9291# 1.15e-19
C183 a_n33_6819# a_18_5680# 1.15e-19
C184 a_n33_n5541# a_18_n5444# 0.0417f
C185 a_18_8152# w_n112_6816# 0.00199f
C186 a_n76_4444# a_n76_3208# 0.00947f
C187 a_n33_n8013# a_n76_n9152# 1.15e-19
C188 a_n76_n7916# a_n33_n9249# 1.15e-19
C189 w_n112_n600# a_n33_n1833# 4.13e-19
C190 a_18_736# a_18_1972# 0.00947f
C191 a_n76_736# a_n33_639# 0.0417f
C192 w_n112_n4308# a_n76_n5444# 0.00199f
C193 a_n76_4444# a_n33_4347# 0.0417f
C194 a_n76_n6680# a_n76_n5444# 0.00947f
C195 a_18_n6680# a_n33_n5541# 1.15e-19
C196 w_n112_n3072# a_n76_n1736# 0.00199f
C197 a_18_8152# a_n76_8152# 0.747f
C198 w_n112_8052# a_18_9388# 0.00199f
C199 w_n112_1872# a_n33_639# 4.13e-19
C200 a_n76_4444# a_n33_5583# 1.15e-19
C201 a_n33_n597# w_n112_n1836# 4.13e-19
C202 a_18_9388# a_n33_9291# 0.0417f
C203 a_n76_3208# a_n33_1875# 1.15e-19
C204 a_n76_n7916# w_n112_n6780# 0.00199f
C205 a_n33_n3069# a_n76_n2972# 0.0417f
C206 a_n33_n9249# a_18_n9152# 0.0417f
C207 a_n76_736# a_n76_n500# 0.00947f
C208 a_18_736# a_n33_n597# 1.15e-19
C209 w_n112_n600# a_18_n1736# 0.00199f
C210 a_18_8152# a_18_6916# 0.00947f
C211 w_n112_n5544# a_n76_n5444# 0.0182f
C212 a_18_4444# w_n112_3108# 0.00199f
C213 a_n33_n5541# a_n33_n6777# 0.0665f
C214 w_n112_n1836# a_n76_n1736# 0.0182f
C215 a_18_n6680# a_18_n5444# 0.00947f
C216 w_n112_n8016# a_n76_n7916# 0.0182f
C217 a_n33_n4305# a_n76_n2972# 1.15e-19
C218 a_18_8152# w_n112_9288# 0.00199f
C219 a_n76_n4208# a_n33_n3069# 1.15e-19
C220 a_18_736# a_n33_639# 0.0417f
C221 a_n76_n6680# w_n112_n5544# 0.00199f
C222 a_n76_3208# w_n112_3108# 0.0182f
C223 a_n76_n7916# w_n112_n9252# 0.00199f
C224 w_n112_4344# a_18_3208# 0.00199f
C225 a_n76_n500# w_n112_n1836# 0.00199f
C226 a_18_9388# a_n76_9388# 0.747f
C227 a_n76_n2972# a_18_n2972# 0.747f
C228 a_n33_4347# w_n112_3108# 4.13e-19
C229 a_n33_n4305# a_n76_n4208# 0.0417f
C230 a_18_1972# a_n33_639# 1.15e-19
C231 a_n33_6819# a_n33_5583# 0.0665f
C232 a_n33_3111# a_18_3208# 0.0417f
C233 a_18_5680# a_18_4444# 0.00947f
C234 a_18_9388# w_n112_9288# 0.0182f
C235 a_n33_n9249# a_n33_n10485# 0.0665f
C236 w_n112_n8016# a_18_n9152# 0.00199f
C237 a_18_n5444# a_n33_n6777# 1.15e-19
C238 a_n33_n9249# a_n76_n9152# 0.0417f
C239 w_n112_4344# a_n76_4444# 0.0182f
C240 a_18_n9152# w_n112_n9252# 0.0182f
C241 w_n112_8052# a_n33_6819# 4.13e-19
C242 a_18_n6680# a_n33_n6777# 0.0417f
C243 a_n76_4444# a_n33_3111# 1.15e-19
C244 w_n112_n3072# a_n76_n2972# 0.0182f
C245 a_n33_n597# a_n33_639# 0.0665f
C246 a_n33_4347# a_18_5680# 1.15e-19
C247 a_n76_n4208# a_18_n4208# 0.747f
C248 a_n33_6819# w_n112_6816# 0.106f
C249 a_n76_n6680# a_n76_n7916# 0.00947f
C250 a_18_n6680# a_n33_n8013# 1.15e-19
C251 a_18_5680# a_n33_5583# 0.0417f
C252 a_n76_1972# a_n33_1875# 0.0417f
C253 a_n33_n10485# a_n76_n10388# 0.0417f
C254 a_18_n500# w_n112_n1836# 0.00199f
C255 a_n33_n597# a_n76_n1736# 1.15e-19
C256 w_n112_1872# a_18_3208# 0.00199f
C257 a_n33_n9249# a_18_n10388# 1.15e-19
C258 a_n76_n9152# a_n76_n10388# 0.00947f
C259 a_n76_n4208# w_n112_n3072# 0.00199f
C260 a_n33_3111# a_n33_1875# 0.0665f
C261 a_n33_6819# a_n76_8152# 1.15e-19
C262 a_18_n9152# w_n112_n10488# 0.00199f
C263 w_n112_n1836# a_n76_n2972# 0.00199f
C264 a_n33_n597# a_n76_n500# 0.0417f
C265 a_18_736# a_18_n500# 0.00947f
C266 w_n112_n8016# a_n76_n9152# 0.00199f
C267 a_18_8152# a_n33_8055# 0.0417f
C268 a_n76_4444# a_n76_5680# 0.00947f
C269 a_n33_n10485# w_n112_n9252# 4.13e-19
C270 a_n33_n1833# a_18_n1736# 0.0417f
C271 a_n33_n8013# a_n33_n6777# 0.0665f
C272 a_18_5680# w_n112_6816# 0.00199f
C273 a_n33_6819# a_18_6916# 0.0417f
C274 a_n76_n9152# w_n112_n9252# 0.0182f
C275 a_18_n6680# a_18_n7916# 0.00947f
C276 a_n76_1972# w_n112_3108# 0.00199f
C277 a_n76_4444# w_n112_5580# 0.00199f
C278 a_n76_n10388# a_18_n10388# 0.747f
C279 a_n76_n500# a_n33_639# 1.15e-19
C280 w_n112_n4308# a_n33_n3069# 4.13e-19
C281 a_n33_4347# a_18_4444# 0.0417f
C282 a_n76_736# a_n33_1875# 1.15e-19
C283 a_n76_n4208# a_n33_n5541# 1.15e-19
C284 a_n33_n4305# a_n76_n5444# 1.15e-19
C285 a_n76_736# w_n112_n600# 0.00199f
C286 a_n33_3111# w_n112_3108# 0.106f
C287 a_18_4444# a_n33_5583# 1.15e-19
C288 a_n76_n500# a_n76_n1736# 0.00947f
C289 w_n112_1872# a_n33_1875# 0.106f
C290 a_18_9388# a_n33_8055# 1.15e-19
C291 a_n76_1972# w_n112_636# 0.00199f
C292 a_n33_4347# a_n76_3208# 1.15e-19
C293 w_n112_n4308# a_n33_n4305# 0.106f
C294 a_n33_n5541# w_n112_n6780# 4.13e-19
C295 a_18_1972# a_18_3208# 0.00947f
C296 a_n33_n10485# w_n112_n10488# 0.106f
C297 a_18_n10388# w_n112_n9252# 0.00199f
C298 w_n112_4344# a_18_5680# 0.00199f
C299 a_n33_n597# a_18_n500# 0.0417f
C300 a_18_n7916# a_n33_n6777# 1.15e-19
C301 a_n76_n9152# w_n112_n10488# 0.00199f
C302 a_18_5680# a_18_6916# 0.00947f
C303 a_n33_4347# a_n33_5583# 0.0665f
C304 w_n112_n4308# a_18_n2972# 0.00199f
C305 a_n33_n1833# a_n33_n3069# 0.0665f
C306 a_n33_6819# a_n76_6916# 0.0417f
C307 a_n33_n8013# a_18_n7916# 0.0417f
C308 a_n33_6819# a_n76_5680# 1.15e-19
C309 a_18_n500# a_n33_639# 1.15e-19
C310 a_18_n10388# VSUBS 0.426f
C311 a_n76_n10388# VSUBS 0.426f
C312 a_n33_n10485# VSUBS 0.192f
C313 a_18_n9152# VSUBS 0.415f
C314 a_n76_n9152# VSUBS 0.415f
C315 a_n33_n9249# VSUBS 0.156f
C316 a_18_n7916# VSUBS 0.415f
C317 a_n76_n7916# VSUBS 0.415f
C318 a_n33_n8013# VSUBS 0.156f
C319 a_18_n6680# VSUBS 0.415f
C320 a_n76_n6680# VSUBS 0.415f
C321 a_n33_n6777# VSUBS 0.156f
C322 a_18_n5444# VSUBS 0.415f
C323 a_n76_n5444# VSUBS 0.415f
C324 a_n33_n5541# VSUBS 0.156f
C325 a_18_n4208# VSUBS 0.415f
C326 a_n76_n4208# VSUBS 0.415f
C327 a_n33_n4305# VSUBS 0.156f
C328 a_18_n2972# VSUBS 0.415f
C329 a_n76_n2972# VSUBS 0.415f
C330 a_n33_n3069# VSUBS 0.156f
C331 a_18_n1736# VSUBS 0.415f
C332 a_n76_n1736# VSUBS 0.415f
C333 a_n33_n1833# VSUBS 0.156f
C334 a_18_n500# VSUBS 0.415f
C335 a_n76_n500# VSUBS 0.415f
C336 a_n33_n597# VSUBS 0.156f
C337 a_18_736# VSUBS 0.415f
C338 a_n76_736# VSUBS 0.415f
C339 a_n33_639# VSUBS 0.156f
C340 a_18_1972# VSUBS 0.415f
C341 a_n76_1972# VSUBS 0.415f
C342 a_n33_1875# VSUBS 0.156f
C343 a_18_3208# VSUBS 0.415f
C344 a_n76_3208# VSUBS 0.415f
C345 a_n33_3111# VSUBS 0.156f
C346 a_18_4444# VSUBS 0.415f
C347 a_n76_4444# VSUBS 0.415f
C348 a_n33_4347# VSUBS 0.156f
C349 a_18_5680# VSUBS 0.415f
C350 a_n76_5680# VSUBS 0.415f
C351 a_n33_5583# VSUBS 0.156f
C352 a_18_6916# VSUBS 0.415f
C353 a_n76_6916# VSUBS 0.415f
C354 a_n33_6819# VSUBS 0.156f
C355 a_18_8152# VSUBS 0.415f
C356 a_n76_8152# VSUBS 0.415f
C357 a_n33_8055# VSUBS 0.156f
C358 a_18_9388# VSUBS 0.426f
C359 a_n76_9388# VSUBS 0.426f
C360 a_n33_9291# VSUBS 0.192f
C361 w_n112_n10488# VSUBS 0.806f
C362 w_n112_n9252# VSUBS 0.806f
C363 w_n112_n8016# VSUBS 0.806f
C364 w_n112_n6780# VSUBS 0.806f
C365 w_n112_n5544# VSUBS 0.806f
C366 w_n112_n4308# VSUBS 0.806f
C367 w_n112_n3072# VSUBS 0.806f
C368 w_n112_n1836# VSUBS 0.806f
C369 w_n112_n600# VSUBS 0.806f
C370 w_n112_636# VSUBS 0.806f
C371 w_n112_1872# VSUBS 0.806f
C372 w_n112_3108# VSUBS 0.806f
C373 w_n112_4344# VSUBS 0.806f
C374 w_n112_5580# VSUBS 0.806f
C375 w_n112_6816# VSUBS 0.806f
C376 w_n112_8052# VSUBS 0.806f
C377 w_n112_9288# VSUBS 0.806f
.ends

.subckt sky130_fd_pr__pfet_01v8_F76D73 a_n1558_11242# a_n1558_n14714# a_n1500_n43239#
+ w_n1594_n3690# a_n1500_n11103# a_n1558_50794# a_1500_n23366# a_n1500_n50655# w_n1594_n56838#
+ w_n1594_n24702# a_1500_n30782# a_n1500_3729# a_n1558_n60446# w_n1594_12378# a_1500_n8534#
+ a_n1558_14950# a_1500_n19658# a_n1500_n14811# a_n1500_n46947# w_n1594_9906# w_n1594_n6162#
+ a_1500_22366# a_n1500_22269# a_n1558_53266# a_n1558_n56738# a_n1558_n24602# a_n1558_21130#
+ a_n1500_n53127# w_n1594_n13578# a_n1558_60682# a_1500_n33254# a_n1500_n60543# w_n1594_n20994#
+ a_1500_n40670# a_1500_18658# a_n1558_49558# a_n1558_17422# w_n1594_22266# a_n1500_n49419#
+ w_n1594_n9870# a_n1500_25977# a_n1558_56974# a_n1500_n56835# a_1500_n29546# a_n1558_n3590#
+ a_1500_n36962# a_n1500_9909# a_n1558_n13478# a_1500_32254# a_n1500_32157# a_n1558_n20894#
+ w_n1594_18558# w_n1594_n23466# a_1500_n43142# w_n1594_n30882# w_n1594_25974# a_n1500_n2451#
+ a_1500_28546# a_1500_n7298# a_n1500_28449# a_n1558_59446# a_n1558_27310# a_n1500_n13575#
+ a_n1500_n59307# w_n1594_32154# w_n1594_n19758# a_1500_35962# a_n1558_n6062# a_n1500_35865#
+ a_1500_n39434# a_n1500_n20991# a_1500_n46850# a_n1558_n23366# a_1500_42142# a_n1500_42045#
+ a_n1558_n30782# w_n1594_n33354# w_n1594_28446# a_1500_n53030# w_n1594_35862# w_n1594_n40770#
+ a_n1558_n9770# w_n1594_18# a_n1558_16186# a_n1500_21# a_n1558_n19658# a_n1500_n16047#
+ a_1500_38434# a_n1500_38337# a_n1500_n55599# a_n1500_n23463# w_n1594_n29646# a_1500_45850#
+ w_n1594_42042# a_n1500_45753# a_n1558_40906# a_1500_n49322# a_n1558_n33254# a_1500_52030#
+ a_n1500_n8631# a_n1558_n40670# a_n1558_19894# w_n1594_38334# w_n1594_n43242# a_n1500_n19755#
+ w_n1594_45750# a_n1558_26074# a_n1558_n29546# a_1500_48322# a_n1500_48225# a_1500_n38198#
+ a_n1558_33490# a_n1558_n36962# a_n1500_n33351# w_n1594_n39534# a_n1500_55641# a_1500_n59210#
+ w_n1594_n46950# a_n1558_n43142# a_n1558_29782# w_n1594_n53130# a_n1500_n29643# w_n1594_48222#
+ a_1500_37198# a_n1558_n39434# a_1500_58210# a_n1500_58113# a_n1500_12381# a_1500_n1118#
+ a_1500_n48086# a_n1558_n46850# w_n1594_n49422# a_n1500_n7395# a_n1558_n53030# w_n1594_37098#
+ a_n1558_39670# a_n1500_n39531# w_n1594_58110# a_1500_n4826# a_1500_47086# a_n1558_10006#
+ a_n1558_n49322# w_n1594_n2454# w_n1594_n38298# a_1500_2590# w_n1594_2490# w_n1594_n59310#
+ a_n1500_6201# a_n1500_18561# a_n1558_13714# a_n1558_2590# a_1500_n25838# a_n1558_n38198#
+ a_1500_5062# a_1500_118# a_n1558_n59210# w_n1594_n48186# w_n1594_n16050# a_1500_n32018#
+ a_n1500_2493# a_1500_24838# a_n1558_5062# a_n1500_n38295# w_n1594_n8634# a_1500_8770#
+ a_n1558_55738# a_n1558_23602# a_n1558_n2354# w_n1594_8670# a_1500_n35726# a_n1558_n48086#
+ a_1500_31018# w_n1594_n58074# w_n1594_24738# a_n1558_8770# a_n1500_n1215# a_n1558_12478#
+ a_n1500_n12339# a_n1500_n48183# a_1500_34726# a_n1500_34629# w_n1594_n25938# a_1500_n45614#
+ a_n1500_8673# w_n1594_n32118# a_n1500_n4923# w_n1594_34626# a_n1558_n8534# w_n1594_n7398#
+ a_n1558_22366# a_n1558_n25838# a_n1500_n22227# a_n1500_n58071# a_1500_44614# a_n1500_44517#
+ a_n1500_n61779# w_n1594_n35826# a_n1500_51933# a_1500_n55502# a_n1558_n32018# a_n1558_18658#
+ w_n1594_n42006# a_n1500_n18519# a_n1500_n25935# w_n1594_44514# w_n1594_51930# a_n1558_32254#
+ a_n1558_n35726# a_n1500_n32115# a_1500_54502# a_n1500_54405# a_1500_n44378# a_1500_n12242#
+ w_n1594_n45714# a_1500_n51794# a_n1500_n3687# a_n1558_28546# a_n1558_n7298# a_n1500_n28407#
+ a_n1558_35962# a_n1500_n35823# w_n1594_54402# a_1500_n15950# a_1500_43378# a_1500_11242#
+ a_n1500_11145# a_n1558_42142# a_n1558_n45614# a_1500_50794# a_n1500_n42003# a_n1500_50697#
+ a_1500_n54266# a_1500_n22130# a_n1500_n6159# w_n1594_n55602# a_1500_n61682# a_n1558_38434#
+ a_n1500_n24699# w_n1594_43278# w_n1594_11142# a_1500_14950# a_n1500_46989# a_n1558_45850#
+ a_n1500_14853# a_1500_n18422# a_n1500_n45711# w_n1594_50694# a_1500_n57974# a_n1500_n9867#
+ w_n1594_n1218# a_1500_53266# a_1500_1354# a_n1500_53169# a_1500_21130# a_n1500_21033#
+ a_n1558_n55502# a_n1558_52030# w_n1594_1254# w_n1594_n12342# w_n1594_n44478# a_1500_60682#
+ a_n1500_60585# w_n1594_14850# w_n1594_n51894# w_n1594_46986# a_1500_49558# a_1500_17422#
+ a_n1558_48322# a_n1500_17325# a_n1500_n34587# a_1500_56974# a_n1558_1354# w_n1594_53166#
+ w_n1594_21030# w_n1594_n4926# a_n1500_56877# a_n1500_24741# a_1500_n3590# a_1500_n28310#
+ w_n1594_60582# w_n1594_4962# a_n1558_n44378# a_n1558_n12242# a_n1558_n51794# w_n1594_17322#
+ w_n1594_n22230# w_n1594_n54366# w_n1594_49458# a_n1500_1257# w_n1594_n61782# w_n1594_56874#
+ a_n1558_37198# a_n1500_n37059# a_1500_59446# a_1500_27310# a_1500_7534# a_n1500_59349#
+ a_n1500_27213# a_1500_n6062# a_1500_n17186# a_n1558_58210# a_n1558_n15950# a_n1500_n44475#
+ a_n1558_n1118# w_n1594_7434# w_n1594_n18522# a_n1500_n51891# a_n1558_n54266# a_1500_n41906#
+ a_n1500_4965# a_n1558_n22130# a_n1558_n61682# w_n1594_59346# w_n1594_27210# a_n1558_7534#
+ a_1500_n9770# w_n1594_30918# a_n1558_n4826# a_1500_16186# a_n1500_16089# a_n1558_47086#
+ a_n1558_n18422# a_n1500_37101# a_n1558_n57974# a_1500_n27074# a_n1500_n54363# a_1500_40906#
+ w_n1594_n28410# a_n1500_40809# a_1500_n34490# a_n1500_7437# w_n1594_16086# a_1500_19894#
+ a_n1500_19797# w_n1594_40806# a_1500_26074# a_1500_6298# a_n1558_n28310# w_n1594_6198#
+ w_n1594_n17286# a_1500_33490# a_n1500_33393# w_n1594_19794# a_n1558_6298# a_1500_29782#
+ a_n1500_29685# a_n1558_24838# w_n1594_33390# a_n1558_n17186# a_n1558_118# a_n1558_31018#
+ w_n1594_n27174# a_n1500_43281# a_n1558_n41906# a_1500_n11006# w_n1594_29682# w_n1594_n34590#
+ a_1500_n50558# a_n1500_n17283# a_1500_39670# a_n1500_39573# a_n1558_34726# a_1500_n14714#
+ a_n1558_n27074# a_1500_10006# a_n1558_n34490# w_n1594_n37062# w_n1594_39570# a_1500_n60446#
+ a_n1500_n27171# a_1500_13714# a_n1500_13617# a_n1500_49461# a_n1558_44614# a_n1500_n30879#
+ a_1500_n56738# a_1500_n24602# w_n1594_n11106# w_n1594_n50658# w_n1594_13614# a_1500_55738#
+ a_1500_23602# a_1500_3826# a_n1500_23505# a_1500_n2354# a_1500_n13478# a_n1558_54502#
+ a_n1500_n40767# w_n1594_3726# w_n1594_n14814# a_n1500_30921# a_1500_n20894# a_n1558_n11006#
+ a_n1558_n50558# w_n1594_n60546# a_n1558_3826# w_n1594_55638# w_n1594_23502# VSUBS
+ a_1500_12478# a_n1558_43378#
X0 a_1500_53266# a_n1500_53169# a_n1558_53266# w_n1594_53166# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1 a_1500_n18422# a_n1500_n18519# a_n1558_n18422# w_n1594_n18522# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X2 a_1500_n45614# a_n1500_n45711# a_n1558_n45614# w_n1594_n45714# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X3 a_1500_n43142# a_n1500_n43239# a_n1558_n43142# w_n1594_n43242# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X4 a_1500_n22130# a_n1500_n22227# a_n1558_n22130# w_n1594_n22230# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X5 a_1500_n3590# a_n1500_n3687# a_n1558_n3590# w_n1594_n3690# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X6 a_1500_35962# a_n1500_35865# a_n1558_35962# w_n1594_35862# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X7 a_1500_33490# a_n1500_33393# a_n1558_33490# w_n1594_33390# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X8 a_1500_60682# a_n1500_60585# a_n1558_60682# w_n1594_60582# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X9 a_1500_12478# a_n1500_12381# a_n1558_12478# w_n1594_12378# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X10 a_1500_38434# a_n1500_38337# a_n1558_38434# w_n1594_38334# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X11 a_1500_6298# a_n1500_6201# a_n1558_6298# w_n1594_6198# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X12 a_1500_n55502# a_n1500_n55599# a_n1558_n55502# w_n1594_n55602# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X13 a_1500_n32018# a_n1500_n32115# a_n1558_n32018# w_n1594_n32118# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X14 a_1500_45850# a_n1500_45753# a_n1558_45850# w_n1594_45750# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X15 a_1500_24838# a_n1500_24741# a_n1558_24838# w_n1594_24738# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X16 a_1500_n38198# a_n1500_n38295# a_n1558_n38198# w_n1594_n38298# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X17 a_1500_22366# a_n1500_22269# a_n1558_22366# w_n1594_22266# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X18 a_1500_48322# a_n1500_48225# a_n1558_48322# w_n1594_48222# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X19 a_1500_n14714# a_n1500_n14811# a_n1558_n14714# w_n1594_n14814# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X20 a_1500_n41906# a_n1500_n42003# a_n1558_n41906# w_n1594_n42006# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X21 a_1500_n12242# a_n1500_n12339# a_n1558_n12242# w_n1594_n12342# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X22 a_1500_34726# a_n1500_34629# a_n1558_34726# w_n1594_34626# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X23 a_1500_32254# a_n1500_32157# a_n1558_32254# w_n1594_32154# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X24 a_1500_n48086# a_n1500_n48183# a_n1558_n48086# w_n1594_n48186# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X25 a_1500_58210# a_n1500_58113# a_n1558_58210# w_n1594_58110# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X26 a_1500_n24602# a_n1500_n24699# a_n1558_n24602# w_n1594_n24702# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X27 a_1500_14950# a_n1500_14853# a_n1558_14950# w_n1594_14850# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X28 a_1500_n8534# a_n1500_n8631# a_n1558_n8534# w_n1594_n8634# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X29 a_1500_n57974# a_n1500_n58071# a_n1558_n57974# w_n1594_n58074# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X30 a_1500_n6062# a_n1500_n6159# a_n1558_n6062# w_n1594_n6162# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X31 a_1500_n34490# a_n1500_n34587# a_n1558_n34490# w_n1594_n34590# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X32 a_1500_17422# a_n1500_17325# a_n1558_17422# w_n1594_17322# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X33 a_1500_44614# a_n1500_44517# a_n1558_44614# w_n1594_44514# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X34 a_1500_42142# a_n1500_42045# a_n1558_42142# w_n1594_42042# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X35 a_1500_8770# a_n1500_8673# a_n1558_8770# w_n1594_8670# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X36 a_1500_n11006# a_n1500_n11103# a_n1558_n11006# w_n1594_n11106# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X37 a_1500_n19658# a_n1500_n19755# a_n1558_n19658# w_n1594_n19758# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X38 a_1500_n46850# a_n1500_n46947# a_n1558_n46850# w_n1594_n46950# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X39 a_1500_n17186# a_n1500_n17283# a_n1558_n17186# w_n1594_n17286# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X40 a_1500_27310# a_n1500_27213# a_n1558_27310# w_n1594_27210# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X41 a_1500_n44378# a_n1500_n44475# a_n1558_n44378# w_n1594_n44478# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X42 a_1500_54502# a_n1500_54405# a_n1558_54502# w_n1594_54402# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X43 a_1500_52030# a_n1500_51933# a_n1558_52030# w_n1594_51930# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X44 a_1500_31018# a_n1500_30921# a_n1558_31018# w_n1594_30918# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X45 a_1500_n4826# a_n1500_n4923# a_n1558_n4826# w_n1594_n4926# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X46 a_1500_37198# a_n1500_37101# a_n1558_37198# w_n1594_37098# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X47 a_1500_n2354# a_n1500_n2451# a_n1558_n2354# w_n1594_n2454# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X48 a_1500_n51794# a_n1500_n51891# a_n1558_n51794# w_n1594_n51894# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X49 a_1500_n29546# a_n1500_n29643# a_n1558_n29546# w_n1594_n29646# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X50 a_1500_13714# a_n1500_13617# a_n1558_13714# w_n1594_13614# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X51 a_1500_n56738# a_n1500_n56835# a_n1558_n56738# w_n1594_n56838# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X52 a_1500_11242# a_n1500_11145# a_n1558_11242# w_n1594_11142# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X53 a_1500_40906# a_n1500_40809# a_n1558_40906# w_n1594_40806# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X54 a_1500_n27074# a_n1500_n27171# a_n1558_n27074# w_n1594_n27174# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X55 a_1500_n54266# a_n1500_n54363# a_n1558_n54266# w_n1594_n54366# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X56 a_1500_19894# a_n1500_19797# a_n1558_19894# w_n1594_19794# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X57 a_1500_2590# a_n1500_2493# a_n1558_2590# w_n1594_2490# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X58 a_1500_n59210# a_n1500_n59307# a_n1558_n59210# w_n1594_n59310# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X59 a_1500_7534# a_n1500_7437# a_n1558_7534# w_n1594_7434# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X60 a_1500_49558# a_n1500_49461# a_n1558_49558# w_n1594_49458# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X61 a_1500_n36962# a_n1500_n37059# a_n1558_n36962# w_n1594_n37062# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X62 a_1500_5062# a_n1500_4965# a_n1558_5062# w_n1594_4962# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X63 a_1500_47086# a_n1500_46989# a_n1558_47086# w_n1594_46986# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X64 a_1500_n15950# a_n1500_n16047# a_n1558_n15950# w_n1594_n16050# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X65 a_1500_n61682# a_n1500_n61779# a_n1558_n61682# w_n1594_n61782# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X66 a_1500_n13478# a_n1500_n13575# a_n1558_n13478# w_n1594_n13578# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X67 a_1500_23602# a_n1500_23505# a_n1558_23602# w_n1594_23502# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X68 a_1500_n40670# a_n1500_n40767# a_n1558_n40670# w_n1594_n40770# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X69 a_1500_n39434# a_n1500_n39531# a_n1558_n39434# w_n1594_n39534# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X70 a_1500_21130# a_n1500_21033# a_n1558_21130# w_n1594_21030# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X71 a_1500_29782# a_n1500_29685# a_n1558_29782# w_n1594_29682# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X72 a_1500_56974# a_n1500_56877# a_n1558_56974# w_n1594_56874# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X73 a_1500_59446# a_n1500_59349# a_n1558_59446# w_n1594_59346# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X74 a_1500_n20894# a_n1500_n20991# a_n1558_n20894# w_n1594_n20994# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X75 a_1500_n25838# a_n1500_n25935# a_n1558_n25838# w_n1594_n25938# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X76 a_1500_n23366# a_n1500_n23463# a_n1558_n23366# w_n1594_n23466# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X77 a_1500_n50558# a_n1500_n50655# a_n1558_n50558# w_n1594_n50658# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X78 a_1500_n49322# a_n1500_n49419# a_n1558_n49322# w_n1594_n49422# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X79 a_1500_n1118# a_n1500_n1215# a_n1558_n1118# w_n1594_n1218# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X80 a_1500_n9770# a_n1500_n9867# a_n1558_n9770# w_n1594_n9870# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X81 a_1500_n28310# a_n1500_n28407# a_n1558_n28310# w_n1594_n28410# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X82 a_1500_n7298# a_n1500_n7395# a_n1558_n7298# w_n1594_n7398# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X83 a_1500_10006# a_n1500_9909# a_n1558_10006# w_n1594_9906# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X84 a_1500_39670# a_n1500_39573# a_n1558_39670# w_n1594_39570# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X85 a_1500_18658# a_n1500_18561# a_n1558_18658# w_n1594_18558# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X86 a_1500_n53030# a_n1500_n53127# a_n1558_n53030# w_n1594_n53130# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X87 a_1500_3826# a_n1500_3729# a_n1558_3826# w_n1594_3726# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X88 a_1500_16186# a_n1500_16089# a_n1558_16186# w_n1594_16086# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X89 a_1500_1354# a_n1500_1257# a_n1558_1354# w_n1594_1254# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X90 a_1500_43378# a_n1500_43281# a_n1558_43378# w_n1594_43278# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X91 a_1500_n30782# a_n1500_n30879# a_n1558_n30782# w_n1594_n30882# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X92 a_1500_118# a_n1500_21# a_n1558_118# w_n1594_18# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X93 a_1500_n35726# a_n1500_n35823# a_n1558_n35726# w_n1594_n35826# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X94 a_1500_n33254# a_n1500_n33351# a_n1558_n33254# w_n1594_n33354# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X95 a_1500_n60446# a_n1500_n60543# a_n1558_n60446# w_n1594_n60546# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X96 a_1500_50794# a_n1500_50697# a_n1558_50794# w_n1594_50694# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X97 a_1500_28546# a_n1500_28449# a_n1558_28546# w_n1594_28446# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X98 a_1500_55738# a_n1500_55641# a_n1558_55738# w_n1594_55638# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X99 a_1500_26074# a_n1500_25977# a_n1558_26074# w_n1594_25974# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
C0 a_n1500_n40767# w_n1594_n39534# 0.0172f
C1 a_1500_n2354# a_1500_n3590# 0.0105f
C2 a_n1500_n3687# a_n1558_n3590# 0.217f
C3 w_n1594_21030# a_n1558_21130# 0.0187f
C4 a_n1500_42045# a_n1500_40809# 3.11f
C5 w_n1594_6198# a_n1500_7437# 0.0172f
C6 w_n1594_n23466# a_n1558_n22130# 0.0023f
C7 a_1500_n19658# a_1500_n20894# 0.0105f
C8 a_n1500_n20991# a_n1558_n20894# 0.217f
C9 a_n1558_n15950# w_n1594_n17286# 0.0023f
C10 w_n1594_n29646# a_1500_n30782# 0.0023f
C11 w_n1594_17322# a_1500_16186# 0.0023f
C12 a_1500_8770# w_n1594_8670# 0.0187f
C13 a_n1558_5062# w_n1594_3726# 0.0023f
C14 w_n1594_19794# a_n1500_19797# 1.65f
C15 a_n1558_n46850# w_n1594_n48186# 0.0023f
C16 a_n1500_48225# a_1500_48322# 0.217f
C17 w_n1594_11142# a_1500_11242# 0.0187f
C18 w_n1594_n8634# a_n1500_n8631# 1.65f
C19 a_1500_52030# a_n1500_51933# 0.217f
C20 w_n1594_n55602# a_n1500_n56835# 0.0172f
C21 a_n1500_22269# w_n1594_23502# 0.0172f
C22 w_n1594_n16050# a_1500_n14714# 0.0023f
C23 a_n1500_n2451# a_n1500_n1215# 3.11f
C24 a_n1500_55641# a_1500_55738# 0.217f
C25 w_n1594_n3690# a_n1558_n3590# 0.0187f
C26 a_n1500_n53127# a_n1500_n54363# 3.11f
C27 a_n1500_27213# w_n1594_27210# 1.65f
C28 a_n1558_34726# w_n1594_34626# 0.0187f
C29 w_n1594_34626# a_1500_33490# 0.0023f
C30 a_n1558_49558# w_n1594_48222# 0.0023f
C31 w_n1594_n34590# a_1500_n35726# 0.0023f
C32 a_n1500_n44475# a_n1500_n45711# 3.11f
C33 w_n1594_n33354# a_n1558_n32018# 0.0023f
C34 w_n1594_40806# a_n1500_40809# 1.65f
C35 w_n1594_n18522# a_1500_n18422# 0.0187f
C36 a_n1558_n57974# a_n1558_n59210# 0.0105f
C37 w_n1594_2490# a_n1500_1257# 0.0172f
C38 w_n1594_25974# a_1500_27310# 0.0023f
C39 w_n1594_n25938# a_n1500_n25935# 1.65f
C40 a_n1500_n11103# a_1500_n11006# 0.217f
C41 a_n1500_4965# a_n1558_5062# 0.217f
C42 w_n1594_14850# a_n1500_16089# 0.0172f
C43 w_n1594_53166# a_n1558_52030# 0.0023f
C44 a_n1558_38434# w_n1594_37098# 0.0023f
C45 a_n1500_n9867# a_n1500_n8631# 3.11f
C46 a_n1558_45850# a_n1558_47086# 0.0105f
C47 w_n1594_29682# a_1500_28546# 0.0023f
C48 w_n1594_n58074# a_1500_n57974# 0.0187f
C49 a_n1500_9909# a_n1500_8673# 3.11f
C50 a_n1558_n38198# w_n1594_n37062# 0.0023f
C51 w_n1594_60582# a_1500_60682# 0.0187f
C52 a_n1558_33490# w_n1594_32154# 0.0023f
C53 w_n1594_n1218# a_1500_n1118# 0.0187f
C54 a_1500_n30782# a_1500_n32018# 0.0105f
C55 a_n1500_n32115# a_n1558_n32018# 0.217f
C56 a_1500_19894# w_n1594_18558# 0.0023f
C57 a_n1500_60585# w_n1594_59346# 0.0172f
C58 a_n1558_n22130# a_n1558_n23366# 0.0105f
C59 a_1500_n44378# w_n1594_n45714# 0.0023f
C60 a_1500_19894# a_1500_18658# 0.0105f
C61 a_n1500_18561# a_n1558_18658# 0.217f
C62 a_n1500_27213# a_n1558_27310# 0.217f
C63 w_n1594_n53130# a_n1558_n54266# 0.0023f
C64 a_1500_28546# a_1500_27310# 0.0105f
C65 a_n1558_n12242# w_n1594_n12342# 0.0187f
C66 a_n1500_n13575# w_n1594_n14814# 0.0172f
C67 a_n1558_n43142# w_n1594_n42006# 0.0023f
C68 w_n1594_n9870# a_1500_n8534# 0.0023f
C69 a_n1500_n39531# w_n1594_n40770# 0.0172f
C70 a_n1500_40809# w_n1594_39570# 0.0172f
C71 a_n1500_44517# a_1500_44614# 0.217f
C72 w_n1594_n20994# a_n1558_n22130# 0.0023f
C73 a_n1500_n61779# a_1500_n61682# 0.217f
C74 w_n1594_n30882# a_1500_n29546# 0.0023f
C75 a_n1500_n16047# a_n1558_n15950# 0.217f
C76 w_n1594_7434# a_1500_7534# 0.0187f
C77 a_1500_n49322# w_n1594_n50658# 0.0023f
C78 a_n1500_21# a_n1500_n1215# 3.11f
C79 a_1500_40906# w_n1594_42042# 0.0023f
C80 a_n1558_n13478# a_n1558_n14714# 0.0105f
C81 w_n1594_53166# a_n1558_53266# 0.0187f
C82 w_n1594_n56838# a_n1500_n55599# 0.0172f
C83 a_n1500_50697# a_n1558_50794# 0.217f
C84 a_1500_52030# a_1500_50794# 0.0105f
C85 a_n1500_n16047# w_n1594_n14814# 0.0172f
C86 a_1500_35962# a_1500_34726# 0.0105f
C87 a_n1558_34726# a_n1558_33490# 0.0105f
C88 a_n1500_34629# a_n1558_34726# 0.217f
C89 w_n1594_n13578# a_n1500_n14811# 0.0172f
C90 a_n1558_n29546# a_n1500_n29643# 0.217f
C91 a_n1500_59349# a_n1500_58113# 3.11f
C92 w_n1594_58110# a_n1500_58113# 1.65f
C93 w_n1594_n35826# a_1500_n34490# 0.0023f
C94 a_1500_45850# w_n1594_44514# 0.0023f
C95 w_n1594_n28410# a_n1558_n28310# 0.0187f
C96 w_n1594_24738# a_1500_23602# 0.0023f
C97 a_n1500_22269# a_n1558_22366# 0.217f
C98 a_1500_23602# a_1500_22366# 0.0105f
C99 w_n1594_n16050# a_n1500_n17283# 0.0172f
C100 a_n1500_n24699# a_n1500_n25935# 3.11f
C101 a_n1558_n36962# a_n1558_n38198# 0.0105f
C102 w_n1594_18# a_n1558_n1118# 0.0023f
C103 w_n1594_n60546# a_n1500_n61779# 0.0172f
C104 a_1500_n40670# w_n1594_n39534# 0.0023f
C105 a_n1500_n3687# a_n1500_n4923# 3.11f
C106 a_n1558_42142# a_n1558_40906# 0.0105f
C107 a_n1558_n36962# w_n1594_n38298# 0.0023f
C108 w_n1594_21030# a_n1500_19797# 0.0172f
C109 w_n1594_6198# a_1500_7534# 0.0023f
C110 a_n1500_n17283# w_n1594_n17286# 1.65f
C111 a_n1500_n20991# a_n1500_n22227# 3.11f
C112 a_n1500_3729# w_n1594_3726# 1.65f
C113 a_n1558_7534# w_n1594_8670# 0.0023f
C114 a_n1558_n49322# a_n1558_n50558# 0.0105f
C115 a_n1500_n48183# w_n1594_n48186# 1.65f
C116 w_n1594_11142# a_n1558_10006# 0.0023f
C117 w_n1594_n55602# a_1500_n56738# 0.0023f
C118 a_1500_22366# w_n1594_23502# 0.0023f
C119 w_n1594_n54366# a_n1558_n53030# 0.0023f
C120 w_n1594_n3690# a_n1500_n4923# 0.0172f
C121 a_n1558_n2354# a_n1558_n1118# 0.0105f
C122 w_n1594_4962# a_n1500_4965# 1.65f
C123 a_n1500_48225# w_n1594_48222# 1.65f
C124 a_n1558_n53030# a_n1558_n54266# 0.0105f
C125 a_n1558_n29546# a_n1558_n30782# 0.0105f
C126 a_n1558_n41906# w_n1594_n43242# 0.0023f
C127 a_n1500_33393# w_n1594_34626# 0.0172f
C128 a_1500_27310# w_n1594_27210# 0.0187f
C129 a_n1558_n44378# a_n1558_n45614# 0.0105f
C130 w_n1594_n33354# a_n1500_n33351# 1.65f
C131 w_n1594_n28410# a_1500_n29546# 0.0023f
C132 w_n1594_40806# a_1500_40906# 0.0187f
C133 w_n1594_40806# a_n1558_39670# 0.0023f
C134 w_n1594_46986# a_n1500_45753# 0.0172f
C135 w_n1594_n30882# a_n1500_n29643# 0.0172f
C136 w_n1594_n18522# a_n1558_n19658# 0.0023f
C137 a_n1500_n59307# a_n1558_n59210# 0.217f
C138 a_1500_n57974# a_1500_n59210# 0.0105f
C139 w_n1594_n25938# a_1500_n25838# 0.0187f
C140 w_n1594_2490# a_1500_1354# 0.0023f
C141 w_n1594_30918# a_n1558_32254# 0.0023f
C142 a_n1500_4965# a_n1500_3729# 3.11f
C143 a_n1500_n40767# a_1500_n40670# 0.217f
C144 w_n1594_14850# a_1500_16186# 0.0023f
C145 a_n1500_37101# w_n1594_37098# 1.65f
C146 a_n1558_n8534# a_n1558_n9770# 0.0105f
C147 a_n1500_n51891# w_n1594_n51894# 1.65f
C148 a_n1558_10006# a_n1558_8770# 0.0105f
C149 w_n1594_n58074# a_n1558_n59210# 0.0023f
C150 a_n1500_32157# w_n1594_32154# 1.65f
C151 a_n1500_n32115# a_n1500_n33351# 3.11f
C152 a_n1558_18658# w_n1594_18558# 0.0187f
C153 w_n1594_n23466# a_1500_n22130# 0.0023f
C154 a_n1558_n45614# w_n1594_n45714# 0.0187f
C155 a_n1500_18561# a_n1500_17325# 3.11f
C156 w_n1594_11142# a_n1500_12381# 0.0172f
C157 a_1500_n13478# w_n1594_n14814# 0.0023f
C158 w_n1594_n19758# a_n1500_n18519# 0.0172f
C159 a_n1500_n56835# a_1500_n56738# 0.217f
C160 a_n1500_n13575# w_n1594_n12342# 0.0172f
C161 w_n1594_n9870# a_n1558_n9770# 0.0187f
C162 w_n1594_n61782# a_n1500_n60543# 0.0172f
C163 a_n1500_n48183# a_1500_n48086# 0.217f
C164 w_n1594_1254# a_n1558_2590# 0.0023f
C165 a_1500_n39434# w_n1594_n40770# 0.0023f
C166 a_1500_40906# w_n1594_39570# 0.0023f
C167 w_n1594_39570# a_n1558_39670# 0.0187f
C168 w_n1594_58110# a_n1500_59349# 0.0172f
C169 w_n1594_n30882# a_n1558_n30782# 0.0187f
C170 a_n1500_n18519# a_1500_n18422# 0.217f
C171 w_n1594_7434# a_n1558_6298# 0.0023f
C172 a_n1500_n16047# a_n1500_n17283# 3.11f
C173 w_n1594_50694# a_n1558_52030# 0.0023f
C174 a_1500_n13478# a_1500_n14714# 0.0105f
C175 a_n1500_n14811# a_n1558_n14714# 0.217f
C176 w_n1594_53166# a_n1500_51933# 0.0172f
C177 a_n1500_50697# a_n1500_49461# 3.11f
C178 w_n1594_n56838# a_1500_n55502# 0.0023f
C179 a_n1500_6201# a_1500_6298# 0.217f
C180 a_1500_34726# a_1500_33490# 0.0105f
C181 a_n1500_33393# a_n1558_33490# 0.217f
C182 a_n1500_34629# a_n1500_33393# 3.11f
C183 a_n1558_33490# a_n1558_32254# 0.0105f
C184 w_n1594_n13578# a_1500_n14714# 0.0023f
C185 w_n1594_n35826# a_n1558_n35726# 0.0187f
C186 a_n1558_44614# w_n1594_44514# 0.0187f
C187 w_n1594_18# a_1500_n1118# 0.0023f
C188 w_n1594_n2454# a_n1558_n1118# 0.0023f
C189 w_n1594_n28410# a_n1500_n29643# 0.0172f
C190 a_n1500_n9867# w_n1594_n11106# 0.0172f
C191 a_n1500_22269# a_n1500_21033# 3.11f
C192 w_n1594_n16050# a_1500_n17186# 0.0023f
C193 a_1500_n36962# a_1500_n38198# 0.0105f
C194 a_n1558_n24602# a_n1558_n25838# 0.0105f
C195 a_n1500_n38295# a_n1558_n38198# 0.217f
C196 a_n1500_n44475# w_n1594_n43242# 0.0172f
C197 w_n1594_n60546# a_1500_n61682# 0.0023f
C198 w_n1594_22266# a_n1558_23602# 0.0023f
C199 w_n1594_n59310# a_n1558_n57974# 0.0023f
C200 a_n1500_40809# a_n1500_39573# 3.11f
C201 a_n1500_40809# a_n1558_40906# 0.217f
C202 a_n1558_n3590# a_n1558_n4826# 0.0105f
C203 a_n1500_n38295# w_n1594_n38298# 1.65f
C204 a_1500_42142# a_1500_40906# 0.0105f
C205 a_n1558_n20894# a_n1558_n22130# 0.0105f
C206 a_1500_n17186# w_n1594_n17286# 0.0187f
C207 w_n1594_6198# a_n1558_6298# 0.0187f
C208 a_n1500_25977# w_n1594_25974# 1.65f
C209 a_1500_3826# w_n1594_3726# 0.0187f
C210 a_n1500_n50655# a_n1558_n50558# 0.217f
C211 a_1500_n48086# w_n1594_n48186# 0.0187f
C212 a_n1500_n37059# a_n1500_n35823# 3.11f
C213 a_n1558_60682# w_n1594_60582# 0.0187f
C214 w_n1594_n20994# a_1500_n22130# 0.0023f
C215 w_n1594_56874# a_n1500_58113# 0.0172f
C216 a_n1500_29685# a_1500_29782# 0.217f
C217 w_n1594_n3690# a_1500_n4826# 0.0023f
C218 w_n1594_n54366# a_n1500_n54363# 1.65f
C219 w_n1594_4962# a_1500_5062# 0.0187f
C220 a_1500_n53030# a_1500_n54266# 0.0105f
C221 a_1500_48322# w_n1594_48222# 0.0187f
C222 a_n1500_n54363# a_n1558_n54266# 0.217f
C223 w_n1594_55638# a_n1500_55641# 1.65f
C224 a_n1500_n43239# w_n1594_n43242# 1.65f
C225 w_n1594_56874# a_n1558_55738# 0.0023f
C226 w_n1594_33390# a_n1558_33490# 0.0187f
C227 w_n1594_33390# a_n1500_34629# 0.0172f
C228 a_1500_21130# a_1500_19894# 0.0105f
C229 a_1500_n44378# a_1500_n45614# 0.0105f
C230 a_n1500_n45711# a_n1558_n45614# 0.217f
C231 w_n1594_n33354# a_1500_n33254# 0.0187f
C232 w_n1594_13614# a_n1558_12478# 0.0023f
C233 w_n1594_59346# a_n1500_58113# 0.0172f
C234 w_n1594_46986# a_1500_45850# 0.0023f
C235 w_n1594_16086# a_n1558_17422# 0.0023f
C236 a_n1500_n59307# a_n1500_n60543# 3.11f
C237 w_n1594_n25938# a_n1558_n27074# 0.0023f
C238 w_n1594_30918# a_n1500_30921# 1.65f
C239 w_n1594_n24702# a_n1500_n23463# 0.0172f
C240 w_n1594_12378# a_n1558_12478# 0.0187f
C241 w_n1594_14850# a_n1558_14950# 0.0187f
C242 a_n1558_5062# a_n1558_3826# 0.0105f
C243 a_n1500_n28407# a_1500_n28310# 0.217f
C244 a_1500_37198# w_n1594_37098# 0.0187f
C245 a_1500_n51794# w_n1594_n51894# 0.0187f
C246 a_n1500_37101# a_1500_37198# 0.217f
C247 a_1500_10006# a_1500_8770# 0.0105f
C248 a_n1500_8673# a_n1558_8770# 0.217f
C249 w_n1594_51930# a_n1558_52030# 0.0187f
C250 a_n1500_n7395# a_1500_n7298# 0.217f
C251 a_1500_32254# w_n1594_32154# 0.0187f
C252 a_n1558_n32018# a_n1558_n33254# 0.0105f
C253 a_n1500_17325# w_n1594_18558# 0.0172f
C254 a_n1558_n15950# a_n1558_n14714# 0.0105f
C255 a_n1500_n46947# w_n1594_n45714# 0.0172f
C256 a_n1558_18658# a_n1558_17422# 0.0105f
C257 a_n1500_24741# a_1500_24838# 0.217f
C258 a_1500_n13478# w_n1594_n12342# 0.0023f
C259 a_n1558_n14714# w_n1594_n14814# 0.0187f
C260 a_n1558_39670# w_n1594_38334# 0.0023f
C261 w_n1594_n19758# a_1500_n18422# 0.0023f
C262 w_n1594_n61782# a_1500_n60446# 0.0023f
C263 w_n1594_n9870# a_n1500_n11103# 0.0172f
C264 w_n1594_1254# a_n1500_1257# 1.65f
C265 a_n1558_n40670# w_n1594_n40770# 0.0187f
C266 w_n1594_39570# a_n1500_38337# 0.0172f
C267 a_n1500_58113# a_1500_58210# 0.217f
C268 w_n1594_n30882# a_n1500_n32115# 0.0172f
C269 w_n1594_50694# a_n1500_50697# 1.65f
C270 a_n1500_56877# a_n1500_55641# 3.11f
C271 a_n1500_11145# w_n1594_9906# 0.0172f
C272 a_n1500_1257# a_1500_1354# 0.217f
C273 w_n1594_13614# a_n1500_14853# 0.0172f
C274 w_n1594_n8634# a_1500_n8534# 0.0187f
C275 a_n1558_50794# a_n1558_49558# 0.0105f
C276 w_n1594_n56838# a_n1558_n56738# 0.0187f
C277 w_n1594_n2454# a_1500_n1118# 0.0023f
C278 w_n1594_n29646# a_n1558_n29546# 0.0187f
C279 a_1500_33490# a_1500_32254# 0.0105f
C280 a_n1500_33393# a_n1500_32157# 3.11f
C281 a_n1500_32157# a_n1558_32254# 0.217f
C282 w_n1594_51930# a_n1558_53266# 0.0023f
C283 w_n1594_35862# a_n1558_37198# 0.0023f
C284 a_n1500_n35823# a_1500_n35726# 0.217f
C285 a_n1500_43281# w_n1594_44514# 0.0172f
C286 w_n1594_n27174# a_n1558_n25838# 0.0023f
C287 a_1500_n9770# w_n1594_n11106# 0.0023f
C288 a_n1500_14853# a_1500_14950# 0.217f
C289 a_n1558_22366# a_n1558_21130# 0.0105f
C290 a_1500_n44378# w_n1594_n43242# 0.0023f
C291 a_1500_n24602# a_1500_n25838# 0.0105f
C292 a_n1500_n25935# a_n1558_n25838# 0.217f
C293 a_n1500_n38295# a_n1500_n39531# 3.11f
C294 a_n1500_25977# w_n1594_27210# 0.0172f
C295 w_n1594_22266# a_n1500_22269# 1.65f
C296 a_n1500_n4923# a_n1558_n4826# 0.217f
C297 w_n1594_46986# a_n1558_48322# 0.0023f
C298 w_n1594_18# a_n1500_1257# 0.0172f
C299 w_n1594_n59310# a_n1500_n59307# 1.65f
C300 a_1500_n3590# a_1500_n4826# 0.0105f
C301 a_1500_n38198# w_n1594_n38298# 0.0187f
C302 a_n1500_39573# a_n1558_39670# 0.217f
C303 a_n1558_40906# a_n1558_39670# 0.0105f
C304 a_n1558_n18422# w_n1594_n17286# 0.0023f
C305 a_n1500_n22227# a_n1558_n22130# 0.217f
C306 w_n1594_n1218# a_n1558_n2354# 0.0023f
C307 w_n1594_59346# a_n1500_59349# 1.65f
C308 w_n1594_50694# a_n1500_51933# 0.0172f
C309 a_n1500_50697# w_n1594_49458# 0.0172f
C310 a_n1558_2590# w_n1594_3726# 0.0023f
C311 a_1500_47086# a_1500_48322# 0.0105f
C312 a_1500_26074# w_n1594_25974# 0.0187f
C313 a_n1558_n49322# w_n1594_n48186# 0.0023f
C314 a_n1500_n45711# w_n1594_n46950# 0.0172f
C315 w_n1594_n54366# a_1500_n54266# 0.0187f
C316 w_n1594_n7398# a_n1500_n6159# 0.0172f
C317 a_n1500_54405# a_1500_54502# 0.217f
C318 w_n1594_4962# a_n1558_3826# 0.0023f
C319 a_n1558_47086# w_n1594_48222# 0.0023f
C320 a_n1500_n54363# a_n1500_n55599# 3.11f
C321 w_n1594_54402# a_n1558_55738# 0.0023f
C322 w_n1594_55638# a_1500_55738# 0.0187f
C323 w_n1594_33390# a_1500_34726# 0.0023f
C324 w_n1594_33390# a_n1500_32157# 0.0172f
C325 a_n1500_19797# a_n1500_18561# 3.11f
C326 a_n1500_n3687# w_n1594_n4926# 0.0172f
C327 a_n1500_n4923# w_n1594_n6162# 0.0172f
C328 a_n1500_n45711# a_n1500_n46947# 3.11f
C329 w_n1594_n33354# a_n1558_n34490# 0.0023f
C330 w_n1594_n32118# a_n1500_n30879# 0.0172f
C331 a_n1558_60682# a_n1558_59446# 0.0105f
C332 w_n1594_16086# a_n1500_16089# 1.65f
C333 a_n1558_n59210# a_n1558_n60446# 0.0105f
C334 a_n1500_n50655# w_n1594_n51894# 0.0172f
C335 w_n1594_30918# a_1500_31018# 0.0187f
C336 a_1500_5062# a_1500_3826# 0.0105f
C337 w_n1594_n24702# a_1500_n23366# 0.0023f
C338 a_n1500_3729# a_n1558_3826# 0.217f
C339 w_n1594_12378# a_n1500_11145# 0.0172f
C340 a_n1500_n12339# a_1500_n12242# 0.217f
C341 w_n1594_14850# a_n1500_13617# 0.0172f
C342 a_n1558_35962# w_n1594_37098# 0.0023f
C343 a_1500_n15950# w_n1594_n14814# 0.0023f
C344 w_n1594_51930# a_n1500_50697# 0.0172f
C345 a_n1500_8673# a_n1500_7437# 3.11f
C346 a_n1558_n53030# w_n1594_n51894# 0.0023f
C347 w_n1594_58110# a_1500_58210# 0.0187f
C348 a_n1558_13714# a_n1558_12478# 0.0105f
C349 a_n1558_31018# w_n1594_32154# 0.0023f
C350 a_n1500_n33351# a_n1558_n33254# 0.217f
C351 a_1500_n32018# a_1500_n33254# 0.0105f
C352 a_1500_17422# w_n1594_18558# 0.0023f
C353 a_1500_n15950# a_1500_n14714# 0.0105f
C354 a_1500_n46850# w_n1594_n45714# 0.0023f
C355 a_n1500_17325# a_n1558_17422# 0.217f
C356 a_1500_18658# a_1500_17422# 0.0105f
C357 a_n1558_44614# w_n1594_43278# 0.0023f
C358 w_n1594_28446# a_n1500_29685# 0.0172f
C359 a_n1500_38337# w_n1594_38334# 1.65f
C360 w_n1594_n19758# a_n1558_n19658# 0.0187f
C361 w_n1594_n9870# a_1500_n11006# 0.0023f
C362 w_n1594_n61782# a_n1558_n61682# 0.0187f
C363 w_n1594_1254# a_1500_1354# 0.0187f
C364 a_n1500_n42003# w_n1594_n40770# 0.0172f
C365 w_n1594_39570# a_1500_38434# 0.0023f
C366 a_n1500_43281# a_1500_43378# 0.217f
C367 w_n1594_n30882# a_1500_n32018# 0.0023f
C368 a_n1558_56974# a_n1558_55738# 0.0105f
C369 w_n1594_50694# a_1500_50794# 0.0187f
C370 a_n1558_n36962# w_n1594_n35826# 0.0023f
C371 a_n1558_n48086# w_n1594_n49422# 0.0023f
C372 a_1500_11242# w_n1594_9906# 0.0023f
C373 a_1500_n49322# a_1500_n50558# 0.0105f
C374 a_1500_n29546# a_n1500_n29643# 0.217f
C375 w_n1594_n8634# a_n1558_n9770# 0.0023f
C376 w_n1594_13614# a_1500_14950# 0.0023f
C377 w_n1594_17322# a_n1558_18658# 0.0023f
C378 a_n1500_49461# a_n1558_49558# 0.217f
C379 a_1500_50794# a_1500_49558# 0.0105f
C380 a_n1500_32157# a_n1500_30921# 3.11f
C381 w_n1594_51930# a_n1500_51933# 1.65f
C382 a_n1558_n50558# w_n1594_n50658# 0.0187f
C383 a_1500_n50558# w_n1594_n49422# 0.0023f
C384 a_n1500_n51891# a_1500_n51794# 0.217f
C385 w_n1594_n34590# a_n1558_n33254# 0.0023f
C386 w_n1594_35862# a_n1500_35865# 1.65f
C387 a_1500_43378# w_n1594_44514# 0.0023f
C388 a_1500_n1118# a_1500_118# 0.0105f
C389 a_n1558_n11006# w_n1594_n11106# 0.0187f
C390 w_n1594_n27174# a_n1500_n27171# 1.65f
C391 a_n1500_21033# a_n1558_21130# 0.217f
C392 a_1500_22366# a_1500_21130# 0.0105f
C393 a_1500_n8534# a_1500_n9770# 0.0105f
C394 a_n1500_n9867# a_n1558_n9770# 0.217f
C395 a_n1558_n38198# a_n1558_n39434# 0.0105f
C396 a_n1500_n25935# a_n1500_n27171# 3.11f
C397 a_1500_26074# w_n1594_27210# 0.0023f
C398 w_n1594_22266# a_1500_22366# 0.0187f
C399 w_n1594_18# a_1500_1354# 0.0023f
C400 w_n1594_46986# a_n1500_46989# 1.65f
C401 a_n1558_n39434# w_n1594_n38298# 0.0023f
C402 w_n1594_n59310# a_1500_n59210# 0.0187f
C403 a_n1500_n4923# a_n1500_n6159# 3.11f
C404 a_n1500_11145# a_1500_11242# 0.217f
C405 a_n1500_39573# a_n1500_38337# 3.11f
C406 w_n1594_19794# a_n1500_18561# 0.0172f
C407 w_n1594_29682# a_n1558_31018# 0.0023f
C408 a_1500_40906# a_1500_39670# 0.0105f
C409 w_n1594_n22230# a_n1500_n23463# 0.0172f
C410 a_n1500_60585# a_1500_60682# 0.217f
C411 a_1500_50794# w_n1594_49458# 0.0023f
C412 a_n1558_24838# w_n1594_25974# 0.0023f
C413 a_1500_n45614# w_n1594_n46950# 0.0023f
C414 w_n1594_n23466# a_n1558_n23366# 0.0187f
C415 w_n1594_n7398# a_1500_n6062# 0.0023f
C416 w_n1594_n54366# a_n1558_n55502# 0.0023f
C417 a_1500_47086# w_n1594_48222# 0.0023f
C418 w_n1594_n53130# a_n1500_n51891# 0.0172f
C419 a_n1558_n35726# w_n1594_n37062# 0.0023f
C420 a_n1500_19797# w_n1594_18558# 0.0172f
C421 a_n1558_n54266# a_n1558_n55502# 0.0105f
C422 w_n1594_55638# a_n1558_54502# 0.0023f
C423 w_n1594_54402# a_n1500_54405# 1.65f
C424 a_n1500_n40767# w_n1594_n42006# 0.0172f
C425 a_1500_n3590# w_n1594_n4926# 0.0023f
C426 a_n1558_19894# a_n1558_18658# 0.0105f
C427 w_n1594_33390# a_1500_32254# 0.0023f
C428 a_n1558_n45614# a_n1558_n46850# 0.0105f
C429 a_1500_n4826# w_n1594_n6162# 0.0023f
C430 a_n1500_45753# a_n1558_45850# 0.217f
C431 w_n1594_n32118# a_1500_n30782# 0.0023f
C432 a_n1558_n15950# a_n1558_n17186# 0.0105f
C433 w_n1594_16086# a_1500_16186# 0.0187f
C434 w_n1594_n20994# a_n1500_n19755# 0.0172f
C435 a_n1500_n60543# a_n1558_n60446# 0.217f
C436 a_n1500_n1215# a_n1558_n1118# 0.217f
C437 a_1500_n59210# a_1500_n60446# 0.0105f
C438 w_n1594_30918# a_n1558_29782# 0.0023f
C439 w_n1594_n24702# a_n1558_n24602# 0.0187f
C440 a_n1500_3729# a_n1500_2493# 3.11f
C441 a_n1500_n42003# a_1500_n41906# 0.217f
C442 w_n1594_14850# a_1500_13714# 0.0023f
C443 w_n1594_12378# a_1500_11242# 0.0023f
C444 a_n1558_43378# w_n1594_42042# 0.0023f
C445 w_n1594_n58074# a_n1500_n56835# 0.0172f
C446 a_n1558_8770# a_n1558_7534# 0.0105f
C447 w_n1594_51930# a_1500_50794# 0.0023f
C448 w_n1594_n56838# a_n1500_n58071# 0.0172f
C449 w_n1594_58110# a_n1558_56974# 0.0023f
C450 a_1500_13714# a_1500_12478# 0.0105f
C451 a_n1500_12381# a_n1558_12478# 0.217f
C452 a_n1500_n33351# a_n1500_n34587# 3.11f
C453 a_n1500_n22227# a_1500_n22130# 0.217f
C454 w_n1594_24738# a_n1558_26074# 0.0023f
C455 a_n1500_n44475# w_n1594_n44478# 1.65f
C456 a_n1500_17325# a_n1500_16089# 3.11f
C457 a_n1500_43281# w_n1594_43278# 1.65f
C458 w_n1594_28446# a_1500_29782# 0.0023f
C459 a_1500_38434# w_n1594_38334# 0.0187f
C460 a_n1500_n23463# a_1500_n23366# 0.217f
C461 w_n1594_n19758# a_n1500_n20991# 0.0172f
C462 a_1500_n41906# w_n1594_n40770# 0.0023f
C463 a_n1500_n49419# a_1500_n49322# 0.217f
C464 w_n1594_6198# a_n1500_4965# 0.0172f
C465 a_n1558_n38198# w_n1594_n39534# 0.0023f
C466 a_n1500_n2451# a_1500_n2354# 0.217f
C467 a_n1500_n19755# a_1500_n19658# 0.217f
C468 w_n1594_60582# a_n1558_59446# 0.0023f
C469 a_n1558_45850# w_n1594_45750# 0.0187f
C470 a_1500_56974# a_1500_55738# 0.0105f
C471 w_n1594_50694# a_n1558_49558# 0.0023f
C472 a_n1500_n50655# a_n1500_n51891# 3.11f
C473 w_n1594_13614# a_n1558_13714# 0.0187f
C474 a_n1558_10006# w_n1594_9906# 0.0187f
C475 a_n1500_9909# w_n1594_8670# 0.0172f
C476 a_n1500_n49419# w_n1594_n49422# 1.65f
C477 w_n1594_17322# a_n1500_17325# 1.65f
C478 a_n1558_n36962# a_n1558_n35726# 0.0105f
C479 a_n1500_49461# a_n1500_48225# 3.11f
C480 w_n1594_56874# a_1500_58210# 0.0023f
C481 a_n1500_n43239# w_n1594_n44478# 0.0172f
C482 w_n1594_n55602# a_n1558_n54266# 0.0023f
C483 a_n1558_24838# w_n1594_23502# 0.0023f
C484 w_n1594_12378# a_n1558_13714# 0.0023f
C485 a_n1558_32254# a_n1558_31018# 0.0105f
C486 w_n1594_n34590# a_n1500_n34587# 1.65f
C487 w_n1594_35862# a_1500_35962# 0.0187f
C488 w_n1594_59346# a_1500_58210# 0.0023f
C489 w_n1594_n18522# a_n1500_n17283# 0.0172f
C490 w_n1594_n27174# a_1500_n27074# 0.0187f
C491 w_n1594_n1218# a_1500_118# 0.0023f
C492 a_n1500_n12339# w_n1594_n11106# 0.0172f
C493 w_n1594_2490# a_n1558_3826# 0.0023f
C494 a_n1500_21033# a_n1500_19797# 3.11f
C495 w_n1594_n16050# a_n1500_n16047# 1.65f
C496 a_n1500_n9867# a_n1500_n11103# 3.11f
C497 a_1500_n38198# a_1500_n39434# 0.0105f
C498 a_n1500_n39531# a_n1558_n39434# 0.217f
C499 a_n1558_n25838# a_n1558_n27074# 0.0105f
C500 a_n1500_n37059# a_1500_n36962# 0.217f
C501 w_n1594_22266# a_n1558_21130# 0.0023f
C502 w_n1594_n59310# a_n1558_n60446# 0.0023f
C503 a_n1558_n4826# a_n1558_n6062# 0.0105f
C504 a_n1558_1354# a_n1558_118# 0.0105f
C505 a_n1558_39670# a_n1558_38434# 0.0105f
C506 w_n1594_19794# a_1500_18658# 0.0023f
C507 a_n1558_59446# a_n1558_58210# 0.0105f
C508 w_n1594_29682# a_n1500_29685# 1.65f
C509 a_n1500_n16047# w_n1594_n17286# 0.0172f
C510 w_n1594_n22230# a_1500_n23366# 0.0023f
C511 a_n1500_n30879# a_1500_n30782# 0.217f
C512 a_n1558_49558# w_n1594_49458# 0.0187f
C513 a_1500_n41906# a_1500_n43142# 0.0105f
C514 a_n1558_n46850# w_n1594_n46950# 0.0187f
C515 w_n1594_n23466# a_n1500_n24699# 0.0172f
C516 w_n1594_n7398# a_n1558_n7298# 0.0187f
C517 a_1500_n1118# a_n1500_n1215# 0.217f
C518 a_n1500_28449# a_1500_28546# 0.217f
C519 w_n1594_n53130# a_1500_n51794# 0.0023f
C520 a_n1500_n55599# a_n1558_n55502# 0.217f
C521 a_1500_n54266# a_1500_n55502# 0.0105f
C522 w_n1594_4962# a_n1500_6201# 0.0172f
C523 a_1500_n40670# w_n1594_n42006# 0.0023f
C524 w_n1594_54402# a_1500_54502# 0.0187f
C525 a_n1558_n4826# w_n1594_n4926# 0.0187f
C526 a_n1558_n6062# w_n1594_n6162# 0.0187f
C527 a_n1500_n46947# a_n1558_n46850# 0.217f
C528 a_1500_n45614# a_1500_n46850# 0.0105f
C529 w_n1594_n32118# a_n1558_n32018# 0.0187f
C530 a_n1500_45753# a_n1500_44517# 3.11f
C531 a_n1500_n17283# a_n1558_n17186# 0.217f
C532 w_n1594_16086# a_n1558_14950# 0.0023f
C533 w_n1594_n20994# a_1500_n19658# 0.0023f
C534 a_n1500_n60543# a_n1500_n61779# 3.11f
C535 a_1500_n15950# a_1500_n17186# 0.0105f
C536 w_n1594_n29646# a_n1558_n28310# 0.0023f
C537 w_n1594_7434# a_n1500_8673# 0.0172f
C538 w_n1594_n24702# a_n1500_n25935# 0.0172f
C539 a_n1558_3826# a_n1558_2590# 0.0105f
C540 a_n1500_42045# w_n1594_42042# 1.65f
C541 w_n1594_n58074# a_1500_n56738# 0.0023f
C542 w_n1594_n2454# a_n1558_n2354# 0.0187f
C543 a_1500_8770# a_1500_7534# 0.0105f
C544 a_n1500_7437# a_n1558_7534# 0.217f
C545 a_n1500_35865# a_1500_35962# 0.217f
C546 w_n1594_n13578# a_n1558_n12242# 0.0023f
C547 w_n1594_n56838# a_1500_n57974# 0.0023f
C548 a_n1500_12381# a_n1500_11145# 3.11f
C549 a_n1558_n33254# a_n1558_n34490# 0.0105f
C550 w_n1594_24738# a_n1500_24741# 1.65f
C551 a_n1500_23505# a_1500_23602# 0.217f
C552 a_n1558_17422# a_n1558_16186# 0.0105f
C553 a_1500_n44378# w_n1594_n44478# 0.0187f
C554 a_1500_43378# w_n1594_43278# 0.0187f
C555 w_n1594_28446# a_n1558_28546# 0.0187f
C556 w_n1594_n19758# a_1500_n20894# 0.0023f
C557 a_n1558_37198# w_n1594_38334# 0.0023f
C558 w_n1594_n22230# a_n1500_n20991# 0.0172f
C559 w_n1594_n60546# a_n1558_n59210# 0.0023f
C560 w_n1594_6198# a_1500_5062# 0.0023f
C561 w_n1594_n9870# a_n1558_n8534# 0.0023f
C562 a_n1500_n39531# w_n1594_n39534# 1.65f
C563 w_n1594_21030# a_n1558_22366# 0.0023f
C564 a_n1500_44517# w_n1594_45750# 0.0172f
C565 w_n1594_n29646# a_1500_n29546# 0.0187f
C566 w_n1594_13614# a_n1500_12381# 0.0172f
C567 a_1500_n49322# w_n1594_n49422# 0.0187f
C568 a_n1500_8673# w_n1594_9906# 0.0172f
C569 a_1500_10006# w_n1594_8670# 0.0023f
C570 a_n1500_60585# a_n1558_60682# 0.217f
C571 w_n1594_17322# a_1500_17422# 0.0187f
C572 w_n1594_19794# a_n1500_21033# 0.0172f
C573 a_1500_n36962# a_1500_n35726# 0.0105f
C574 a_n1558_49558# a_n1558_48322# 0.0105f
C575 w_n1594_56874# a_n1558_56974# 0.0187f
C576 w_n1594_55638# a_n1500_56877# 0.0172f
C577 w_n1594_11142# a_1500_12478# 0.0023f
C578 w_n1594_n8634# a_n1500_n7395# 0.0172f
C579 a_n1500_23505# w_n1594_23502# 1.65f
C580 w_n1594_n55602# a_n1500_n55599# 1.65f
C581 a_n1558_52030# a_n1558_53266# 0.0105f
C582 w_n1594_12378# a_n1500_12381# 1.65f
C583 w_n1594_n3690# a_n1558_n2354# 0.0023f
C584 a_n1500_30921# a_n1558_31018# 0.217f
C585 a_1500_32254# a_1500_31018# 0.0105f
C586 a_n1500_28449# w_n1594_27210# 0.0172f
C587 a_n1558_35962# w_n1594_34626# 0.0023f
C588 a_n1500_59349# a_1500_59446# 0.217f
C589 w_n1594_n34590# a_1500_n34490# 0.0187f
C590 w_n1594_58110# a_1500_59446# 0.0023f
C591 w_n1594_35862# a_n1558_34726# 0.0023f
C592 w_n1594_40806# a_n1500_42045# 0.0172f
C593 w_n1594_n18522# a_1500_n17186# 0.0023f
C594 w_n1594_1254# a_1500_118# 0.0023f
C595 a_1500_n12242# w_n1594_n11106# 0.0023f
C596 w_n1594_n27174# a_n1558_n28310# 0.0023f
C597 a_n1500_n58071# a_1500_n57974# 0.217f
C598 a_n1558_21130# a_n1558_19894# 0.0105f
C599 a_n1500_13617# a_1500_13714# 0.217f
C600 w_n1594_2490# a_n1500_2493# 1.65f
C601 w_n1594_n25938# a_n1500_n24699# 0.0172f
C602 a_n1558_n9770# a_n1558_n11006# 0.0105f
C603 a_n1500_n39531# a_n1500_n40767# 3.11f
C604 a_1500_n25838# a_1500_n27074# 0.0105f
C605 a_n1500_n27171# a_n1558_n27074# 0.217f
C606 a_n1500_n6159# a_n1558_n6062# 0.217f
C607 a_1500_1354# a_1500_118# 0.0105f
C608 w_n1594_29682# a_1500_29782# 0.0187f
C609 a_n1500_21# a_n1558_118# 0.217f
C610 a_1500_n4826# a_1500_n6062# 0.0105f
C611 a_n1500_38337# a_n1558_38434# 0.217f
C612 a_n1558_n36962# w_n1594_n37062# 0.0187f
C613 a_n1500_n37059# w_n1594_n38298# 0.0172f
C614 a_1500_39670# a_1500_38434# 0.0105f
C615 a_n1500_48225# w_n1594_49458# 0.0172f
C616 a_n1500_n43239# a_n1500_n44475# 3.11f
C617 a_n1500_n48183# w_n1594_n46950# 0.0172f
C618 w_n1594_n23466# a_1500_n24602# 0.0023f
C619 a_n1500_25977# a_n1558_26074# 0.217f
C620 a_n1500_53169# a_1500_53266# 0.217f
C621 w_n1594_n7398# a_n1500_n8631# 0.0172f
C622 w_n1594_n53130# a_n1558_n53030# 0.0187f
C623 a_n1500_n55599# a_n1500_n56835# 3.11f
C624 w_n1594_4962# a_1500_6298# 0.0023f
C625 w_n1594_54402# a_n1558_53266# 0.0023f
C626 a_n1558_n11006# w_n1594_n12342# 0.0023f
C627 a_n1558_n41906# w_n1594_n42006# 0.0187f
C628 w_n1594_n1218# a_n1500_n1215# 1.65f
C629 a_n1500_n6159# w_n1594_n4926# 0.0172f
C630 a_n1500_n7395# w_n1594_n6162# 0.0172f
C631 a_n1500_n46947# a_n1500_n48183# 3.11f
C632 a_n1558_45850# a_n1558_44614# 0.0105f
C633 w_n1594_n32118# a_n1500_n33351# 0.0172f
C634 w_n1594_n20994# a_n1558_n20894# 0.0187f
C635 a_n1500_n17283# a_n1500_n18519# 3.11f
C636 a_n1558_n60446# a_n1558_n61682# 0.0105f
C637 w_n1594_n29646# a_n1500_n29643# 1.65f
C638 w_n1594_7434# a_1500_8770# 0.0023f
C639 w_n1594_18# a_1500_118# 0.0187f
C640 w_n1594_n24702# a_1500_n25838# 0.0023f
C641 a_n1500_2493# a_n1558_2590# 0.217f
C642 a_1500_3826# a_1500_2590# 0.0105f
C643 a_1500_42142# w_n1594_42042# 0.0187f
C644 a_n1500_n13575# a_1500_n13478# 0.217f
C645 w_n1594_53166# a_n1558_54502# 0.0023f
C646 w_n1594_n2454# a_n1500_n3687# 0.0172f
C647 a_n1500_7437# a_n1500_6201# 3.11f
C648 a_n1500_n51891# w_n1594_n50658# 0.0172f
C649 w_n1594_n13578# a_n1500_n13575# 1.65f
C650 a_n1500_n34587# a_n1558_n34490# 0.217f
C651 a_1500_n33254# a_1500_n34490# 0.0105f
C652 w_n1594_n28410# a_n1558_n27074# 0.0023f
C653 w_n1594_24738# a_1500_24838# 0.0187f
C654 a_n1500_16089# a_n1558_16186# 0.217f
C655 a_1500_17422# a_1500_16186# 0.0105f
C656 a_n1558_n45614# w_n1594_n44478# 0.0023f
C657 a_n1558_42142# w_n1594_43278# 0.0023f
C658 w_n1594_28446# a_n1500_27213# 0.0172f
C659 w_n1594_n22230# a_1500_n20894# 0.0023f
C660 w_n1594_n60546# a_n1500_n60543# 1.65f
C661 a_1500_n39434# w_n1594_n39534# 0.0187f
C662 a_n1500_42045# a_1500_42142# 0.217f
C663 w_n1594_21030# a_n1500_21033# 1.65f
C664 w_n1594_n23466# a_n1500_n22227# 0.0172f
C665 w_n1594_n29646# a_n1558_n30782# 0.0023f
C666 a_1500_44614# w_n1594_45750# 0.0023f
C667 a_1500_8770# w_n1594_9906# 0.0023f
C668 a_n1500_4965# w_n1594_3726# 0.0172f
C669 a_n1558_8770# w_n1594_8670# 0.0187f
C670 a_n1500_n46947# w_n1594_n48186# 0.0172f
C671 w_n1594_19794# a_1500_21130# 0.0023f
C672 w_n1594_17322# a_n1558_16186# 0.0023f
C673 w_n1594_11142# a_n1558_11242# 0.0187f
C674 a_n1500_48225# a_n1558_48322# 0.217f
C675 a_1500_49558# a_1500_48322# 0.0105f
C676 w_n1594_55638# a_1500_56974# 0.0023f
C677 w_n1594_n8634# a_1500_n7298# 0.0023f
C678 a_n1558_52030# a_n1500_51933# 0.217f
C679 a_1500_52030# a_1500_53266# 0.0105f
C680 w_n1594_n16050# a_n1558_n14714# 0.0023f
C681 w_n1594_n55602# a_1500_n55502# 0.0187f
C682 a_1500_23602# w_n1594_23502# 0.0187f
C683 w_n1594_n3690# a_n1500_n3687# 1.65f
C684 a_n1500_55641# a_n1558_55738# 0.217f
C685 a_n1500_30921# a_n1500_29685# 3.11f
C686 a_n1500_n53127# a_1500_n53030# 0.217f
C687 w_n1594_34626# a_n1558_33490# 0.0023f
C688 a_n1500_49461# w_n1594_48222# 0.0172f
C689 a_n1500_34629# w_n1594_34626# 1.65f
C690 a_1500_28546# w_n1594_27210# 0.0023f
C691 w_n1594_n34590# a_n1558_n35726# 0.0023f
C692 a_n1500_n44475# a_1500_n44378# 0.217f
C693 w_n1594_n33354# a_n1500_n32115# 0.0172f
C694 w_n1594_n18522# a_n1558_n18422# 0.0187f
C695 w_n1594_40806# a_1500_42142# 0.0023f
C696 a_n1500_19797# a_n1558_19894# 0.217f
C697 w_n1594_25974# a_n1558_27310# 0.0023f
C698 w_n1594_n25938# a_1500_n24602# 0.0023f
C699 w_n1594_2490# a_1500_2590# 0.0187f
C700 a_1500_n9770# a_1500_n11006# 0.0105f
C701 a_n1500_n11103# a_n1558_n11006# 0.217f
C702 a_n1500_n27171# a_n1500_n28407# 3.11f
C703 a_n1558_n39434# a_n1558_n40670# 0.0105f
C704 a_n1500_38337# w_n1594_37098# 0.0172f
C705 a_1500_n8534# a_n1500_n8631# 0.217f
C706 w_n1594_n58074# a_n1558_n57974# 0.0187f
C707 w_n1594_29682# a_n1558_28546# 0.0023f
C708 a_n1500_n6159# a_n1500_n7395# 3.11f
C709 a_n1500_9909# a_1500_10006# 0.217f
C710 a_n1500_38337# a_n1500_37101# 3.11f
C711 a_n1500_n38295# w_n1594_n37062# 0.0172f
C712 a_1500_48322# w_n1594_49458# 0.0023f
C713 a_n1558_n43142# a_n1558_n44378# 0.0105f
C714 a_n1500_60585# w_n1594_60582# 1.65f
C715 a_1500_n48086# w_n1594_n46950# 0.0023f
C716 a_n1558_n44378# w_n1594_n45714# 0.0023f
C717 a_n1500_25977# a_n1500_24741# 3.11f
C718 w_n1594_n53130# a_n1500_n54363# 0.0172f
C719 a_n1558_n55502# a_n1558_n56738# 0.0105f
C720 a_n1500_n12339# w_n1594_n12342# 1.65f
C721 a_n1500_n43239# w_n1594_n42006# 0.0172f
C722 a_1500_n6062# w_n1594_n4926# 0.0023f
C723 a_n1500_56877# a_1500_56974# 0.217f
C724 a_1500_n7298# w_n1594_n6162# 0.0023f
C725 a_n1558_n46850# a_n1558_n48086# 0.0105f
C726 a_1500_45850# a_1500_44614# 0.0105f
C727 a_n1500_44517# a_n1558_44614# 0.217f
C728 w_n1594_59346# a_1500_59446# 0.0187f
C729 w_n1594_n32118# a_1500_n33254# 0.0023f
C730 a_n1558_n17186# a_n1558_n18422# 0.0105f
C731 a_n1500_n61779# a_n1558_n61682# 0.217f
C732 w_n1594_n20994# a_n1500_n22227# 0.0172f
C733 a_1500_n60446# a_1500_n61682# 0.0105f
C734 w_n1594_7434# a_n1558_7534# 0.0187f
C735 a_n1558_n49322# w_n1594_n50658# 0.0023f
C736 a_n1500_2493# a_n1500_1257# 3.11f
C737 a_n1558_40906# w_n1594_42042# 0.0023f
C738 w_n1594_53166# a_n1500_53169# 1.65f
C739 w_n1594_n2454# a_1500_n3590# 0.0023f
C740 a_n1558_7534# a_n1558_6298# 0.0105f
C741 a_n1558_47086# w_n1594_45750# 0.0023f
C742 a_1500_n51794# w_n1594_n50658# 0.0023f
C743 w_n1594_n13578# a_1500_n13478# 0.0187f
C744 w_n1594_n35826# a_n1558_n34490# 0.0023f
C745 a_n1500_n34587# a_n1500_n35823# 3.11f
C746 a_n1558_45850# w_n1594_44514# 0.0023f
C747 w_n1594_n28410# a_n1500_n28407# 1.65f
C748 w_n1594_24738# a_n1558_23602# 0.0023f
C749 a_n1500_16089# a_n1500_14853# 3.11f
C750 w_n1594_n16050# a_1500_n15950# 0.0187f
C751 w_n1594_28446# a_1500_27310# 0.0023f
C752 a_n1500_n24699# a_1500_n24602# 0.217f
C753 w_n1594_n22230# a_n1558_n22130# 0.0187f
C754 w_n1594_18# a_n1500_n1215# 0.0172f
C755 w_n1594_n60546# a_1500_n60446# 0.0187f
C756 a_n1558_n40670# w_n1594_n39534# 0.0023f
C757 a_n1500_n3687# a_1500_n3590# 0.217f
C758 w_n1594_21030# a_1500_21130# 0.0187f
C759 a_1500_59446# a_1500_58210# 0.0105f
C760 w_n1594_6198# a_n1558_7534# 0.0023f
C761 a_n1500_n20991# a_1500_n20894# 0.217f
C762 a_1500_n15950# w_n1594_n17286# 0.0023f
C763 a_1500_5062# w_n1594_3726# 0.0023f
C764 a_n1500_7437# w_n1594_8670# 0.0172f
C765 a_1500_n46850# w_n1594_n48186# 0.0023f
C766 w_n1594_19794# a_n1558_19894# 0.0187f
C767 w_n1594_n8634# a_n1558_n8534# 0.0187f
C768 w_n1594_11142# a_n1500_9909# 0.0172f
C769 a_n1500_48225# a_n1500_46989# 3.11f
C770 a_n1500_50697# a_n1500_51933# 3.11f
C771 a_n1558_22366# w_n1594_23502# 0.0023f
C772 w_n1594_n55602# a_n1558_n56738# 0.0023f
C773 w_n1594_n54366# a_n1500_n53127# 0.0172f
C774 a_n1500_55641# a_n1500_54405# 3.11f
C775 w_n1594_n3690# a_1500_n3590# 0.0187f
C776 a_n1558_31018# a_n1558_29782# 0.0105f
C777 a_1500_49558# w_n1594_48222# 0.0023f
C778 a_1500_34726# w_n1594_34626# 0.0187f
C779 a_n1558_27310# w_n1594_27210# 0.0187f
C780 a_n1558_n50558# a_n1558_n51794# 0.0105f
C781 a_n1500_n42003# w_n1594_n43242# 0.0172f
C782 w_n1594_n33354# a_1500_n32018# 0.0023f
C783 w_n1594_40806# a_n1500_39573# 0.0172f
C784 w_n1594_40806# a_n1558_40906# 0.0187f
C785 w_n1594_n18522# a_n1500_n19755# 0.0172f
C786 w_n1594_30918# a_n1500_32157# 0.0172f
C787 w_n1594_n25938# a_n1558_n25838# 0.0187f
C788 w_n1594_2490# a_n1558_1354# 0.0023f
C789 w_n1594_14850# a_n1558_16186# 0.0023f
C790 a_n1500_4965# a_1500_5062# 0.217f
C791 a_1500_n39434# a_1500_n40670# 0.0105f
C792 a_n1500_n11103# a_n1500_n12339# 3.11f
C793 w_n1594_53166# a_1500_52030# 0.0023f
C794 a_n1500_n40767# a_n1558_n40670# 0.217f
C795 a_n1558_n27074# a_n1558_n28310# 0.0105f
C796 a_1500_38434# w_n1594_37098# 0.0023f
C797 w_n1594_n58074# a_n1500_n59307# 0.0172f
C798 a_1500_n50558# w_n1594_n51894# 0.0023f
C799 a_n1558_n6062# a_n1558_n7298# 0.0105f
C800 a_1500_n38198# w_n1594_n37062# 0.0023f
C801 a_n1558_38434# a_n1558_37198# 0.0105f
C802 a_1500_33490# w_n1594_32154# 0.0023f
C803 w_n1594_59346# a_1500_60682# 0.0023f
C804 a_n1500_n32115# a_1500_n32018# 0.217f
C805 a_n1500_18561# w_n1594_18558# 1.65f
C806 a_n1500_n45711# w_n1594_n45714# 1.65f
C807 a_n1558_26074# a_n1558_24838# 0.0105f
C808 a_n1500_18561# a_1500_18658# 0.217f
C809 a_n1500_27213# a_1500_27310# 0.217f
C810 w_n1594_n53130# a_1500_n54266# 0.0023f
C811 a_n1500_n56835# a_n1558_n56738# 0.217f
C812 a_1500_n55502# a_1500_n56738# 0.0105f
C813 a_1500_n12242# w_n1594_n12342# 0.0187f
C814 a_n1558_n13478# w_n1594_n14814# 0.0023f
C815 w_n1594_n9870# a_n1500_n9867# 1.65f
C816 a_n1500_n48183# a_n1558_n48086# 0.217f
C817 a_n1558_n39434# w_n1594_n40770# 0.0023f
C818 a_1500_n46850# a_1500_n48086# 0.0105f
C819 w_n1594_1254# a_n1500_2493# 0.0172f
C820 w_n1594_39570# a_n1500_39573# 1.65f
C821 a_n1558_40906# w_n1594_39570# 0.0023f
C822 a_n1500_44517# a_n1500_43281# 3.11f
C823 a_1500_n17186# a_1500_n18422# 0.0105f
C824 a_n1500_n18519# a_n1558_n18422# 0.217f
C825 w_n1594_n30882# a_n1500_n30879# 1.65f
C826 a_n1500_n16047# a_1500_n15950# 0.217f
C827 w_n1594_7434# a_n1500_6201# 0.0172f
C828 a_n1500_n50655# w_n1594_n50658# 1.65f
C829 a_n1558_2590# a_n1558_1354# 0.0105f
C830 w_n1594_53166# a_1500_53266# 0.0187f
C831 w_n1594_n56838# a_n1558_n55502# 0.0023f
C832 a_n1500_50697# a_1500_50794# 0.217f
C833 a_1500_47086# w_n1594_45750# 0.0023f
C834 a_1500_7534# a_1500_6298# 0.0105f
C835 a_n1500_6201# a_n1558_6298# 0.217f
C836 a_n1500_34629# a_1500_34726# 0.217f
C837 w_n1594_n13578# a_n1558_n14714# 0.0023f
C838 w_n1594_n35826# a_n1500_n35823# 1.65f
C839 a_n1500_44517# w_n1594_44514# 1.65f
C840 a_n1558_n34490# a_n1558_n35726# 0.0105f
C841 w_n1594_n2454# a_n1500_n1215# 0.0172f
C842 w_n1594_n28410# a_1500_n28310# 0.0187f
C843 a_n1558_16186# a_n1558_14950# 0.0105f
C844 a_n1500_22269# a_1500_22366# 0.217f
C845 w_n1594_n16050# a_n1558_n17186# 0.0023f
C846 a_1500_n43142# w_n1594_n43242# 0.0187f
C847 w_n1594_22266# a_n1500_23505# 0.0172f
C848 w_n1594_n60546# a_n1558_n61682# 0.0023f
C849 w_n1594_n59310# a_n1500_n58071# 0.0172f
C850 w_n1594_21030# a_n1558_19894# 0.0023f
C851 a_1500_n36962# w_n1594_n38298# 0.0023f
C852 a_n1558_n17186# w_n1594_n17286# 0.0187f
C853 w_n1594_6198# a_n1500_6201# 1.65f
C854 a_n1500_n37059# w_n1594_n35826# 0.0172f
C855 a_1500_7534# w_n1594_8670# 0.0023f
C856 a_n1558_3826# w_n1594_3726# 0.0187f
C857 a_n1558_n48086# w_n1594_n48186# 0.0187f
C858 w_n1594_n7398# a_1500_n8534# 0.0023f
C859 w_n1594_11142# a_1500_10006# 0.0023f
C860 a_n1558_48322# a_n1558_47086# 0.0105f
C861 w_n1594_n54366# a_1500_n53030# 0.0023f
C862 a_n1558_55738# a_n1558_54502# 0.0105f
C863 a_1500_31018# a_1500_29782# 0.0105f
C864 w_n1594_n3690# a_n1558_n4826# 0.0023f
C865 a_n1500_29685# a_n1558_29782# 0.217f
C866 w_n1594_4962# a_n1558_5062# 0.0187f
C867 a_n1558_48322# w_n1594_48222# 0.0187f
C868 a_1500_n41906# w_n1594_n43242# 0.0023f
C869 w_n1594_56874# a_n1500_55641# 0.0172f
C870 a_n1558_n50558# w_n1594_n49422# 0.0023f
C871 w_n1594_n33354# a_n1558_n33254# 0.0187f
C872 w_n1594_40806# a_1500_39670# 0.0023f
C873 w_n1594_46986# a_n1558_45850# 0.0023f
C874 w_n1594_n18522# a_1500_n19658# 0.0023f
C875 w_n1594_16086# a_n1500_17325# 0.0172f
C876 a_n1500_n59307# a_1500_n59210# 0.217f
C877 w_n1594_30918# a_1500_32254# 0.0023f
C878 w_n1594_n25938# a_n1500_n27171# 0.0172f
C879 w_n1594_14850# a_n1500_14853# 1.65f
C880 a_n1558_n11006# a_n1558_n12242# 0.0105f
C881 a_n1500_n40767# a_n1500_n42003# 3.11f
C882 a_n1558_37198# w_n1594_37098# 0.0187f
C883 a_1500_n27074# a_1500_n28310# 0.0105f
C884 a_n1500_n28407# a_n1558_n28310# 0.217f
C885 a_1500_47086# a_1500_45850# 0.0105f
C886 w_n1594_n58074# a_1500_n59210# 0.0023f
C887 a_n1500_n7395# a_n1558_n7298# 0.217f
C888 a_n1500_37101# a_n1558_37198# 0.217f
C889 a_1500_38434# a_1500_37198# 0.0105f
C890 a_n1558_n51794# w_n1594_n51894# 0.0187f
C891 a_1500_n6062# a_1500_n7298# 0.0105f
C892 w_n1594_n22230# a_1500_n22130# 0.0187f
C893 a_n1558_32254# w_n1594_32154# 0.0187f
C894 a_n1500_33393# w_n1594_32154# 0.0172f
C895 a_1500_18658# w_n1594_18558# 0.0187f
C896 a_1500_n45614# w_n1594_n45714# 0.0187f
C897 a_n1500_24741# a_n1558_24838# 0.217f
C898 a_1500_26074# a_1500_24838# 0.0105f
C899 a_n1558_n13478# w_n1594_n12342# 0.0023f
C900 a_n1500_n14811# w_n1594_n14814# 1.65f
C901 a_n1500_39573# w_n1594_38334# 0.0172f
C902 w_n1594_n19758# a_n1558_n18422# 0.0023f
C903 w_n1594_n61782# a_n1558_n60446# 0.0023f
C904 w_n1594_n9870# a_1500_n9770# 0.0187f
C905 w_n1594_1254# a_1500_2590# 0.0023f
C906 a_n1500_n40767# w_n1594_n40770# 1.65f
C907 a_n1500_n48183# a_n1500_n49419# 3.11f
C908 a_n1500_58113# a_n1558_58210# 0.217f
C909 w_n1594_39570# a_1500_39670# 0.0187f
C910 a_n1558_44614# a_n1558_43378# 0.0105f
C911 w_n1594_n30882# a_1500_n30782# 0.0187f
C912 a_n1500_n18519# a_n1500_n19755# 3.11f
C913 w_n1594_7434# a_1500_6298# 0.0023f
C914 w_n1594_50694# a_1500_52030# 0.0023f
C915 a_n1500_n14811# a_1500_n14714# 0.217f
C916 a_n1500_1257# a_n1558_1354# 0.217f
C917 a_1500_2590# a_1500_1354# 0.0105f
C918 w_n1594_n56838# a_n1500_n56835# 1.65f
C919 a_n1500_33393# a_1500_33490# 0.217f
C920 w_n1594_51930# a_n1500_53169# 0.0172f
C921 w_n1594_n35826# a_1500_n35726# 0.0187f
C922 w_n1594_35862# a_n1500_37101# 0.0172f
C923 a_1500_n34490# a_1500_n35726# 0.0105f
C924 a_n1500_n35823# a_n1558_n35726# 0.217f
C925 a_1500_44614# w_n1594_44514# 0.0187f
C926 a_n1558_n9770# w_n1594_n11106# 0.0023f
C927 w_n1594_n27174# a_n1500_n25935# 0.0172f
C928 a_1500_16186# a_1500_14950# 0.0105f
C929 a_n1500_14853# a_n1558_14950# 0.217f
C930 a_n1500_n38295# a_1500_n38198# 0.217f
C931 a_n1558_n44378# w_n1594_n43242# 0.0023f
C932 a_1500_n22130# a_1500_n23366# 0.0105f
C933 w_n1594_22266# a_1500_23602# 0.0023f
C934 a_n1558_118# a_n1558_n1118# 0.0105f
C935 w_n1594_46986# a_n1500_48225# 0.0172f
C936 w_n1594_n59310# a_1500_n57974# 0.0023f
C937 a_n1558_12478# a_n1558_11242# 0.0105f
C938 a_n1500_40809# a_1500_40906# 0.217f
C939 a_n1558_n38198# w_n1594_n38298# 0.0187f
C940 a_1500_n1118# a_1500_n2354# 0.0105f
C941 w_n1594_6198# a_1500_6298# 0.0187f
C942 a_n1500_n18519# w_n1594_n17286# 0.0172f
C943 w_n1594_60582# a_n1500_59349# 0.0172f
C944 w_n1594_n1218# a_n1500_n2451# 0.0172f
C945 a_n1558_26074# w_n1594_25974# 0.0187f
C946 a_n1500_2493# w_n1594_3726# 0.0172f
C947 a_n1500_n49419# w_n1594_n48186# 0.0172f
C948 a_n1558_60682# w_n1594_59346# 0.0023f
C949 a_n1500_46989# a_n1558_47086# 0.217f
C950 a_1500_55738# a_1500_54502# 0.0105f
C951 w_n1594_n54366# a_n1558_n54266# 0.0187f
C952 a_n1500_29685# a_n1500_28449# 3.11f
C953 a_n1500_54405# a_n1558_54502# 0.217f
C954 w_n1594_4962# a_n1500_3729# 0.0172f
C955 a_n1500_n54363# a_1500_n54266# 0.217f
C956 a_n1500_46989# w_n1594_48222# 0.0172f
C957 w_n1594_56874# a_1500_55738# 0.0023f
C958 a_n1558_n43142# w_n1594_n43242# 0.0187f
C959 w_n1594_54402# a_n1500_55641# 0.0172f
C960 w_n1594_55638# a_n1558_55738# 0.0187f
C961 w_n1594_33390# a_n1558_34726# 0.0023f
C962 w_n1594_33390# a_1500_33490# 0.0187f
C963 a_n1500_19797# a_1500_19894# 0.217f
C964 a_n1500_n56835# a_n1500_n58071# 3.11f
C965 a_n1500_n45711# a_1500_n45614# 0.217f
C966 w_n1594_n33354# a_n1500_n34587# 0.0172f
C967 w_n1594_13614# a_1500_12478# 0.0023f
C968 w_n1594_16086# a_1500_17422# 0.0023f
C969 w_n1594_n25938# a_1500_n27074# 0.0023f
C970 w_n1594_30918# a_n1558_31018# 0.0187f
C971 w_n1594_n24702# a_n1558_n23366# 0.0023f
C972 a_1500_n11006# a_1500_n12242# 0.0105f
C973 w_n1594_12378# a_1500_12478# 0.0187f
C974 a_n1500_n12339# a_n1558_n12242# 0.217f
C975 a_n1558_n40670# a_n1558_n41906# 0.0105f
C976 w_n1594_14850# a_1500_14950# 0.0187f
C977 a_n1500_25977# a_n1500_27213# 3.11f
C978 a_n1500_n28407# a_n1500_n29643# 3.11f
C979 a_n1500_35865# w_n1594_37098# 0.0172f
C980 a_n1558_n15950# w_n1594_n14814# 0.0023f
C981 a_n1500_8673# a_1500_8770# 0.217f
C982 w_n1594_51930# a_1500_52030# 0.0187f
C983 a_n1500_n7395# a_n1500_n8631# 3.11f
C984 a_n1500_n53127# w_n1594_n51894# 0.0172f
C985 a_n1500_37101# a_n1500_35865# 3.11f
C986 w_n1594_58110# a_n1558_58210# 0.0187f
C987 a_n1500_30921# w_n1594_32154# 0.0172f
C988 a_n1558_17422# w_n1594_18558# 0.0023f
C989 a_n1558_n46850# w_n1594_n45714# 0.0023f
C990 a_n1500_24741# a_n1500_23505# 3.11f
C991 a_n1500_44517# w_n1594_43278# 0.0172f
C992 w_n1594_n19758# a_n1500_n19755# 1.65f
C993 a_1500_39670# w_n1594_38334# 0.0023f
C994 a_1500_n14714# w_n1594_n14814# 0.0187f
C995 w_n1594_n9870# a_n1558_n11006# 0.0023f
C996 w_n1594_n61782# a_n1500_n61779# 1.65f
C997 a_n1558_n48086# a_n1558_n49322# 0.0105f
C998 w_n1594_n1218# a_n1500_21# 0.0172f
C999 a_1500_n40670# w_n1594_n40770# 0.0187f
C1000 w_n1594_1254# a_n1558_1354# 0.0187f
C1001 a_n1500_58113# a_n1500_56877# 3.11f
C1002 w_n1594_39570# a_n1558_38434# 0.0023f
C1003 a_n1500_43281# a_n1558_43378# 0.217f
C1004 a_1500_44614# a_1500_43378# 0.0105f
C1005 w_n1594_n30882# a_n1558_n32018# 0.0023f
C1006 a_n1558_n18422# a_n1558_n19658# 0.0105f
C1007 w_n1594_50694# a_n1558_50794# 0.0187f
C1008 a_n1500_1257# a_n1500_21# 3.11f
C1009 a_n1500_n48183# w_n1594_n49422# 0.0172f
C1010 a_n1558_11242# w_n1594_9906# 0.0023f
C1011 w_n1594_n8634# a_n1500_n9867# 0.0172f
C1012 w_n1594_13614# a_n1558_14950# 0.0023f
C1013 w_n1594_17322# a_n1500_18561# 0.0172f
C1014 a_1500_n29546# a_1500_n28310# 0.0105f
C1015 w_n1594_n56838# a_1500_n56738# 0.0187f
C1016 a_n1500_32157# a_1500_32254# 0.217f
C1017 a_1500_n50558# a_1500_n51794# 0.0105f
C1018 w_n1594_51930# a_1500_53266# 0.0023f
C1019 a_n1500_n51891# a_n1558_n51794# 0.217f
C1020 w_n1594_n34590# a_n1500_n33351# 0.0172f
C1021 w_n1594_35862# a_1500_37198# 0.0023f
C1022 a_n1558_43378# w_n1594_44514# 0.0023f
C1023 w_n1594_n27174# a_1500_n25838# 0.0023f
C1024 a_n1500_n11103# w_n1594_n11106# 1.65f
C1025 a_n1500_14853# a_n1500_13617# 3.11f
C1026 a_n1500_n25935# a_1500_n25838# 0.217f
C1027 w_n1594_22266# a_n1558_22366# 0.0187f
C1028 a_n1558_26074# w_n1594_27210# 0.0023f
C1029 w_n1594_n59310# a_n1558_n59210# 0.0187f
C1030 a_1500_12478# a_1500_11242# 0.0105f
C1031 w_n1594_46986# a_1500_48322# 0.0023f
C1032 a_n1500_n4923# a_1500_n4826# 0.217f
C1033 w_n1594_18# a_n1558_1354# 0.0023f
C1034 a_n1500_11145# a_n1558_11242# 0.217f
C1035 a_1500_n18422# w_n1594_n17286# 0.0023f
C1036 w_n1594_19794# a_1500_19894# 0.0187f
C1037 a_n1500_39573# a_1500_39670# 0.217f
C1038 w_n1594_29682# a_n1500_30921# 0.0172f
C1039 a_n1500_n39531# w_n1594_n38298# 0.0172f
C1040 w_n1594_n1218# a_1500_n2354# 0.0023f
C1041 a_1500_47086# a_n1500_46989# 0.217f
C1042 a_1500_2590# w_n1594_3726# 0.0023f
C1043 a_n1558_50794# w_n1594_49458# 0.0023f
C1044 a_n1500_24741# w_n1594_25974# 0.0172f
C1045 a_1500_n49322# w_n1594_n48186# 0.0023f
C1046 w_n1594_n23466# a_n1500_n23463# 1.65f
C1047 a_n1558_n45614# w_n1594_n46950# 0.0023f
C1048 w_n1594_n7398# a_n1558_n6062# 0.0023f
C1049 w_n1594_n54366# a_n1500_n55599# 0.0172f
C1050 a_n1500_54405# a_n1500_53169# 3.11f
C1051 a_n1558_29782# a_n1558_28546# 0.0105f
C1052 w_n1594_4962# a_1500_3826# 0.0023f
C1053 a_n1500_n35823# w_n1594_n37062# 0.0172f
C1054 w_n1594_54402# a_1500_55738# 0.0023f
C1055 w_n1594_55638# a_n1500_54405# 0.0172f
C1056 w_n1594_33390# a_n1500_33393# 1.65f
C1057 a_n1558_n3590# w_n1594_n4926# 0.0023f
C1058 w_n1594_33390# a_n1558_32254# 0.0023f
C1059 a_n1558_n4826# w_n1594_n6162# 0.0023f
C1060 a_n1558_n56738# a_n1558_n57974# 0.0105f
C1061 a_1500_60682# a_1500_59446# 0.0105f
C1062 a_n1500_59349# a_n1558_59446# 0.217f
C1063 w_n1594_58110# a_n1558_59446# 0.0023f
C1064 w_n1594_n33354# a_1500_n34490# 0.0023f
C1065 w_n1594_n32118# a_n1558_n30782# 0.0023f
C1066 w_n1594_16086# a_n1558_16186# 0.0187f
C1067 w_n1594_30918# a_n1500_29685# 0.0172f
C1068 a_n1500_3729# a_1500_3826# 0.217f
C1069 w_n1594_n24702# a_n1500_n24699# 1.65f
C1070 a_n1500_n42003# a_n1558_n41906# 0.217f
C1071 w_n1594_14850# a_n1558_13714# 0.0023f
C1072 a_n1500_43281# w_n1594_42042# 0.0172f
C1073 w_n1594_12378# a_n1558_11242# 0.0023f
C1074 a_n1500_n12339# a_n1500_n13575# 3.11f
C1075 a_1500_n40670# a_1500_n41906# 0.0105f
C1076 a_n1558_26074# a_n1558_27310# 0.0105f
C1077 a_1500_35962# w_n1594_37098# 0.0023f
C1078 a_n1500_4965# a_n1500_6201# 3.11f
C1079 a_n1558_n8534# a_n1558_n7298# 0.0105f
C1080 w_n1594_51930# a_n1558_50794# 0.0023f
C1081 a_1500_n53030# w_n1594_n51894# 0.0023f
C1082 a_n1558_37198# a_n1558_35962# 0.0105f
C1083 a_n1500_n37059# w_n1594_n37062# 1.65f
C1084 w_n1594_58110# a_n1500_56877# 0.0172f
C1085 a_1500_31018# w_n1594_32154# 0.0023f
C1086 a_n1500_n33351# a_1500_n33254# 0.217f
C1087 w_n1594_24738# a_n1500_25977# 0.0172f
C1088 a_1500_n20894# a_1500_n22130# 0.0105f
C1089 a_1500_n43142# w_n1594_n44478# 0.0023f
C1090 a_n1558_24838# a_n1558_23602# 0.0105f
C1091 a_n1500_17325# a_1500_17422# 0.217f
C1092 a_1500_44614# w_n1594_43278# 0.0023f
C1093 w_n1594_28446# a_n1558_29782# 0.0023f
C1094 a_n1500_n23463# a_n1558_n23366# 0.217f
C1095 w_n1594_n19758# a_1500_n19658# 0.0187f
C1096 a_n1558_38434# w_n1594_38334# 0.0187f
C1097 w_n1594_n61782# a_1500_n61682# 0.0187f
C1098 w_n1594_1254# a_n1500_21# 0.0172f
C1099 a_n1558_n41906# w_n1594_n40770# 0.0023f
C1100 a_1500_n48086# a_1500_n49322# 0.0105f
C1101 a_n1500_n49419# a_n1558_n49322# 0.217f
C1102 a_n1500_n38295# w_n1594_n39534# 0.0172f
C1103 a_n1500_43281# a_n1500_42045# 3.11f
C1104 a_n1500_n2451# a_n1558_n2354# 0.217f
C1105 a_1500_n18422# a_1500_n19658# 0.0105f
C1106 a_n1500_n19755# a_n1558_n19658# 0.217f
C1107 a_n1500_45753# w_n1594_45750# 1.65f
C1108 a_1500_n36962# w_n1594_n35826# 0.0023f
C1109 w_n1594_50694# a_n1500_49461# 0.0172f
C1110 a_1500_n48086# w_n1594_n49422# 0.0023f
C1111 a_n1500_n50655# a_1500_n50558# 0.217f
C1112 a_n1500_9909# w_n1594_9906# 1.65f
C1113 a_n1500_n30879# a_n1500_n29643# 3.11f
C1114 w_n1594_17322# a_1500_18658# 0.0023f
C1115 w_n1594_n8634# a_1500_n9770# 0.0023f
C1116 w_n1594_13614# a_n1500_13617# 1.65f
C1117 a_n1500_49461# a_1500_49558# 0.217f
C1118 w_n1594_56874# a_n1558_58210# 0.0023f
C1119 a_n1500_24741# w_n1594_23502# 0.0172f
C1120 w_n1594_n55602# a_n1500_n54363# 0.0172f
C1121 w_n1594_12378# a_n1500_13617# 0.0172f
C1122 a_n1500_n51891# a_n1500_n53127# 3.11f
C1123 w_n1594_n34590# a_1500_n33254# 0.0023f
C1124 w_n1594_59346# a_n1558_58210# 0.0023f
C1125 w_n1594_35862# a_n1558_35962# 0.0187f
C1126 w_n1594_n27174# a_n1558_n27074# 0.0187f
C1127 a_1500_n11006# w_n1594_n11106# 0.0187f
C1128 w_n1594_n1218# a_n1558_118# 0.0023f
C1129 w_n1594_2490# a_n1500_3729# 0.0172f
C1130 a_n1558_14950# a_n1558_13714# 0.0105f
C1131 a_n1500_21033# a_1500_21130# 0.217f
C1132 a_n1500_n9867# a_1500_n9770# 0.217f
C1133 w_n1594_21030# a_1500_19894# 0.0023f
C1134 a_n1500_n37059# a_n1558_n36962# 0.217f
C1135 w_n1594_22266# a_n1500_21033# 0.0172f
C1136 w_n1594_n59310# a_n1500_n60543# 0.0172f
C1137 w_n1594_46986# a_n1558_47086# 0.0187f
C1138 w_n1594_18# a_n1500_21# 1.65f
C1139 a_1500_n39434# w_n1594_n38298# 0.0023f
C1140 a_n1500_11145# a_n1500_9909# 3.11f
C1141 w_n1594_29682# a_1500_31018# 0.0023f
C1142 w_n1594_19794# a_n1558_18658# 0.0023f
C1143 w_n1594_n22230# a_n1558_n23366# 0.0023f
C1144 a_n1500_n30879# a_n1558_n30782# 0.217f
C1145 a_n1500_49461# w_n1594_49458# 1.65f
C1146 a_1500_24838# w_n1594_25974# 0.0023f
C1147 a_1500_n29546# a_1500_n30782# 0.0105f
C1148 a_n1500_n46947# w_n1594_n46950# 1.65f
C1149 w_n1594_n23466# a_1500_n23366# 0.0187f
C1150 w_n1594_n7398# a_n1500_n7395# 1.65f
C1151 a_n1500_28449# a_n1558_28546# 0.217f
C1152 w_n1594_n54366# a_1500_n55502# 0.0023f
C1153 a_1500_29782# a_1500_28546# 0.0105f
C1154 a_n1558_54502# a_n1558_53266# 0.0105f
C1155 a_1500_n35726# w_n1594_n37062# 0.0023f
C1156 w_n1594_n53130# a_n1558_n51794# 0.0023f
C1157 a_n1558_19894# w_n1594_18558# 0.0023f
C1158 w_n1594_55638# a_1500_54502# 0.0023f
C1159 a_n1558_n40670# w_n1594_n42006# 0.0023f
C1160 w_n1594_54402# a_n1558_54502# 0.0187f
C1161 a_n1500_n4923# w_n1594_n4926# 1.65f
C1162 a_1500_n56738# a_1500_n57974# 0.0105f
C1163 a_n1500_n6159# w_n1594_n6162# 1.65f
C1164 a_n1500_45753# a_1500_45850# 0.217f
C1165 w_n1594_n32118# a_n1500_n32115# 1.65f
C1166 a_n1500_n60543# a_1500_n60446# 0.217f
C1167 w_n1594_16086# a_n1500_14853# 0.0172f
C1168 w_n1594_n20994# a_n1558_n19658# 0.0023f
C1169 w_n1594_n29646# a_n1500_n28407# 0.0172f
C1170 w_n1594_30918# a_1500_29782# 0.0023f
C1171 w_n1594_n24702# a_1500_n24602# 0.0187f
C1172 a_1500_43378# w_n1594_42042# 0.0023f
C1173 a_n1500_n42003# a_n1500_n43239# 3.11f
C1174 a_n1558_n12242# a_n1558_n13478# 0.0105f
C1175 a_1500_26074# a_1500_27310# 0.0105f
C1176 a_n1558_5062# a_n1558_6298# 0.0105f
C1177 w_n1594_n30882# a_n1558_n29546# 0.0023f
C1178 w_n1594_n58074# a_n1558_n56738# 0.0023f
C1179 a_n1558_n8534# a_n1500_n8631# 0.217f
C1180 w_n1594_n2454# a_n1500_n2451# 1.65f
C1181 a_n1500_35865# a_n1558_35962# 0.217f
C1182 a_1500_37198# a_1500_35962# 0.0105f
C1183 w_n1594_n13578# a_n1500_n12339# 0.0172f
C1184 w_n1594_n56838# a_n1558_n57974# 0.0023f
C1185 w_n1594_58110# a_1500_56974# 0.0023f
C1186 a_n1500_12381# a_1500_12478# 0.217f
C1187 w_n1594_24738# a_1500_26074# 0.0023f
C1188 a_n1500_23505# a_n1558_23602# 0.217f
C1189 a_1500_24838# a_1500_23602# 0.0105f
C1190 a_n1558_n44378# w_n1594_n44478# 0.0187f
C1191 a_n1558_43378# w_n1594_43278# 0.0187f
C1192 w_n1594_28446# a_n1500_28449# 1.65f
C1193 w_n1594_n19758# a_n1558_n20894# 0.0023f
C1194 a_n1500_n23463# a_n1500_n24699# 3.11f
C1195 a_n1500_37101# w_n1594_38334# 0.0172f
C1196 w_n1594_6198# a_n1558_5062# 0.0023f
C1197 w_n1594_n60546# a_n1500_n59307# 0.0172f
C1198 a_n1500_n49419# a_n1500_n50655# 3.11f
C1199 a_1500_n38198# w_n1594_n39534# 0.0023f
C1200 w_n1594_n9870# a_n1500_n8631# 0.0172f
C1201 a_n1558_43378# a_n1558_42142# 0.0105f
C1202 a_n1500_n2451# a_n1500_n3687# 3.11f
C1203 w_n1594_21030# a_n1500_22269# 0.0172f
C1204 a_n1500_n19755# a_n1500_n20991# 3.11f
C1205 a_1500_45850# w_n1594_45750# 0.0187f
C1206 w_n1594_59346# a_n1558_59446# 0.0187f
C1207 w_n1594_50694# a_1500_49558# 0.0023f
C1208 w_n1594_13614# a_1500_13714# 0.0187f
C1209 a_n1558_n49322# w_n1594_n49422# 0.0187f
C1210 a_1500_10006# w_n1594_9906# 0.0187f
C1211 a_n1558_10006# w_n1594_8670# 0.0023f
C1212 w_n1594_17322# a_n1558_17422# 0.0187f
C1213 w_n1594_56874# a_n1500_56877# 1.65f
C1214 w_n1594_11142# a_n1558_12478# 0.0023f
C1215 a_1500_24838# w_n1594_23502# 0.0023f
C1216 a_n1558_n43142# w_n1594_n44478# 0.0023f
C1217 w_n1594_n55602# a_1500_n54266# 0.0023f
C1218 w_n1594_n3690# a_n1500_n2451# 0.0172f
C1219 w_n1594_12378# a_1500_13714# 0.0023f
C1220 a_n1558_n51794# a_n1558_n53030# 0.0105f
C1221 a_n1500_35865# w_n1594_34626# 0.0172f
C1222 w_n1594_n34590# a_n1558_n34490# 0.0187f
C1223 w_n1594_35862# a_n1500_34629# 0.0172f
C1224 w_n1594_n18522# a_n1558_n17186# 0.0023f
C1225 w_n1594_n27174# a_n1500_n28407# 0.0172f
C1226 a_n1500_n58071# a_n1558_n57974# 0.217f
C1227 a_n1558_n12242# w_n1594_n11106# 0.0023f
C1228 w_n1594_1254# a_n1558_118# 0.0023f
C1229 a_1500_14950# a_1500_13714# 0.0105f
C1230 a_n1500_13617# a_n1558_13714# 0.217f
C1231 w_n1594_2490# a_1500_3826# 0.0023f
C1232 a_n1500_n39531# a_1500_n39434# 0.217f
C1233 w_n1594_n28410# a_n1558_n29546# 0.0023f
C1234 a_n1500_n37059# a_n1500_n38295# 3.11f
C1235 w_n1594_46986# a_1500_47086# 0.0187f
C1236 w_n1594_22266# a_1500_21130# 0.0023f
C1237 w_n1594_n59310# a_1500_n60446# 0.0023f
C1238 a_n1558_11242# a_n1558_10006# 0.0105f
C1239 w_n1594_29682# a_n1558_29782# 0.0187f
C1240 a_1500_49558# w_n1594_49458# 0.0187f
C1241 a_n1500_n43239# a_1500_n43142# 0.217f
C1242 a_n1500_n30879# a_n1500_n32115# 3.11f
C1243 a_1500_n46850# w_n1594_n46950# 0.0187f
C1244 w_n1594_n23466# a_n1558_n24602# 0.0023f
C1245 a_n1500_53169# a_n1558_53266# 0.217f
C1246 w_n1594_n7398# a_1500_n7298# 0.0187f
C1247 a_1500_54502# a_1500_53266# 0.0105f
C1248 a_n1500_28449# a_n1500_27213# 3.11f
C1249 w_n1594_n53130# a_n1500_n53127# 1.65f
C1250 a_n1500_n55599# a_1500_n55502# 0.217f
C1251 w_n1594_4962# a_n1558_6298# 0.0023f
C1252 a_n1500_n42003# w_n1594_n42006# 1.65f
C1253 a_n1500_n11103# w_n1594_n12342# 0.0172f
C1254 w_n1594_54402# a_n1500_53169# 0.0172f
C1255 a_1500_n4826# w_n1594_n4926# 0.0187f
C1256 a_n1558_58210# a_n1558_56974# 0.0105f
C1257 a_n1500_n46947# a_1500_n46850# 0.217f
C1258 a_1500_n6062# w_n1594_n6162# 0.0187f
C1259 w_n1594_n32118# a_1500_n32018# 0.0187f
C1260 a_n1500_n17283# a_1500_n17186# 0.217f
C1261 w_n1594_16086# a_1500_14950# 0.0023f
C1262 w_n1594_n20994# a_n1500_n20991# 1.65f
C1263 w_n1594_n29646# a_1500_n28310# 0.0023f
C1264 w_n1594_7434# a_n1558_8770# 0.0023f
C1265 w_n1594_18# a_n1558_118# 0.0187f
C1266 w_n1594_n24702# a_n1558_n25838# 0.0023f
C1267 a_n1558_42142# w_n1594_42042# 0.0187f
C1268 a_n1558_n41906# a_n1558_n43142# 0.0105f
C1269 a_1500_n12242# a_1500_n13478# 0.0105f
C1270 a_n1500_n13575# a_n1558_n13478# 0.217f
C1271 w_n1594_53166# a_n1500_54405# 0.0172f
C1272 a_1500_5062# a_1500_6298# 0.0105f
C1273 w_n1594_n2454# a_1500_n2354# 0.0187f
C1274 a_n1500_7437# a_1500_7534# 0.217f
C1275 a_n1558_n50558# w_n1594_n51894# 0.0023f
C1276 a_1500_n50558# w_n1594_n50658# 0.0187f
C1277 a_n1500_35865# a_n1500_34629# 3.11f
C1278 w_n1594_n13578# a_1500_n12242# 0.0023f
C1279 w_n1594_n28410# a_n1500_n27171# 0.0172f
C1280 w_n1594_24738# a_n1558_24838# 0.0187f
C1281 a_n1500_23505# a_n1500_22269# 3.11f
C1282 a_n1500_n45711# w_n1594_n44478# 0.0172f
C1283 a_n1500_42045# w_n1594_43278# 0.0172f
C1284 w_n1594_28446# a_1500_28546# 0.0187f
C1285 a_1500_37198# w_n1594_38334# 0.0023f
C1286 w_n1594_n22230# a_n1558_n20894# 0.0023f
C1287 a_n1558_n23366# a_n1558_n24602# 0.0105f
C1288 w_n1594_n60546# a_1500_n59210# 0.0023f
C1289 a_n1558_n39434# w_n1594_n39534# 0.0187f
C1290 a_1500_43378# a_1500_42142# 0.0105f
C1291 w_n1594_21030# a_1500_22366# 0.0023f
C1292 a_n1500_42045# a_n1558_42142# 0.217f
C1293 a_n1558_n2354# a_n1558_n3590# 0.0105f
C1294 a_n1558_n19658# a_n1558_n20894# 0.0105f
C1295 a_n1558_44614# w_n1594_45750# 0.0023f
C1296 w_n1594_n29646# a_n1500_n30879# 0.0172f
C1297 a_n1500_60585# a_n1500_59349# 3.11f
C1298 a_n1500_n50655# w_n1594_n49422# 0.0172f
C1299 a_n1558_8770# w_n1594_9906# 0.0023f
C1300 a_n1500_8673# w_n1594_8670# 1.65f
C1301 w_n1594_19794# a_n1558_21130# 0.0023f
C1302 w_n1594_17322# a_n1500_16089# 0.0172f
C1303 w_n1594_56874# a_1500_56974# 0.0187f
C1304 w_n1594_55638# a_n1558_56974# 0.0023f
C1305 w_n1594_11142# a_n1500_11145# 1.65f
C1306 w_n1594_n8634# a_n1558_n7298# 0.0023f
C1307 w_n1594_n16050# a_n1500_n14811# 0.0172f
C1308 w_n1594_n55602# a_n1558_n55502# 0.0187f
C1309 a_n1558_23602# w_n1594_23502# 0.0187f
C1310 w_n1594_n3690# a_1500_n2354# 0.0023f
C1311 a_n1500_30921# a_1500_31018# 0.217f
C1312 a_1500_n51794# a_1500_n53030# 0.0105f
C1313 a_n1500_n53127# a_n1558_n53030# 0.217f
C1314 a_1500_35962# w_n1594_34626# 0.0023f
C1315 a_n1558_28546# w_n1594_27210# 0.0023f
C1316 a_1500_n43142# a_1500_n44378# 0.0105f
C1317 a_n1500_n44475# a_n1558_n44378# 0.217f
C1318 w_n1594_n34590# a_n1500_n35823# 0.0172f
C1319 w_n1594_35862# a_1500_34726# 0.0023f
C1320 w_n1594_n18522# a_n1500_n18519# 1.65f
C1321 w_n1594_40806# a_n1558_42142# 0.0023f
C1322 w_n1594_n27174# a_1500_n28310# 0.0023f
C1323 a_n1500_n58071# a_n1500_n59307# 3.11f
C1324 w_n1594_n25938# a_n1558_n24602# 0.0023f
C1325 w_n1594_2490# a_n1558_2590# 0.0187f
C1326 a_n1500_13617# a_n1500_12381# 3.11f
C1327 w_n1594_25974# a_n1500_27213# 0.0172f
C1328 a_n1500_n27171# a_1500_n27074# 0.217f
C1329 a_1500_n43142# w_n1594_n42006# 0.0023f
C1330 a_1500_n8534# a_1500_n7298# 0.0105f
C1331 a_n1500_45753# a_n1500_46989# 3.11f
C1332 a_n1500_21# a_1500_118# 0.217f
C1333 w_n1594_n58074# a_n1500_n58071# 1.65f
C1334 a_1500_11242# a_1500_10006# 0.0105f
C1335 a_n1500_9909# a_n1558_10006# 0.217f
C1336 a_n1500_n6159# a_1500_n6062# 0.217f
C1337 w_n1594_29682# a_n1500_28449# 0.0172f
C1338 a_n1500_38337# a_1500_38434# 0.217f
C1339 a_1500_n36962# w_n1594_n37062# 0.0187f
C1340 a_n1558_n30782# a_n1558_n32018# 0.0105f
C1341 a_n1558_48322# w_n1594_49458# 0.0023f
C1342 a_n1500_n22227# a_n1500_n23463# 3.11f
C1343 a_n1558_n48086# w_n1594_n46950# 0.0023f
C1344 a_n1500_n44475# w_n1594_n45714# 0.0172f
C1345 w_n1594_n7398# a_n1558_n8534# 0.0023f
C1346 a_n1500_25977# a_1500_26074# 0.217f
C1347 a_n1500_53169# a_n1500_51933# 3.11f
C1348 w_n1594_n53130# a_1500_n53030# 0.0187f
C1349 a_n1558_28546# a_n1558_27310# 0.0105f
C1350 a_1500_n11006# w_n1594_n12342# 0.0023f
C1351 w_n1594_54402# a_1500_53266# 0.0023f
C1352 w_n1594_n1218# a_n1558_n1118# 0.0187f
C1353 a_1500_n41906# w_n1594_n42006# 0.0187f
C1354 a_n1500_56877# a_n1558_56974# 0.217f
C1355 a_1500_58210# a_1500_56974# 0.0105f
C1356 a_n1558_n6062# w_n1594_n4926# 0.0023f
C1357 a_n1558_n7298# w_n1594_n6162# 0.0023f
C1358 w_n1594_n32118# a_n1558_n33254# 0.0023f
C1359 w_n1594_60582# a_1500_59446# 0.0023f
C1360 w_n1594_n20994# a_1500_n20894# 0.0187f
C1361 w_n1594_7434# a_n1500_7437# 1.65f
C1362 a_n1500_n49419# w_n1594_n50658# 0.0172f
C1363 a_n1500_2493# a_1500_2590# 0.217f
C1364 a_n1500_40809# w_n1594_42042# 0.0172f
C1365 a_n1500_n43239# a_n1558_n43142# 0.217f
C1366 a_n1500_n13575# a_n1500_n14811# 3.11f
C1367 w_n1594_53166# a_1500_54502# 0.0023f
C1368 a_n1558_52030# a_n1558_50794# 0.0105f
C1369 w_n1594_n2454# a_n1558_n3590# 0.0023f
C1370 a_n1558_35962# a_n1558_34726# 0.0105f
C1371 a_n1500_46989# w_n1594_45750# 0.0172f
C1372 a_n1558_n51794# w_n1594_n50658# 0.0023f
C1373 w_n1594_n13578# a_n1558_n13478# 0.0187f
C1374 a_n1558_n29546# a_n1558_n28310# 0.0105f
C1375 w_n1594_n35826# a_n1500_n34587# 0.0172f
C1376 a_n1500_n34587# a_1500_n34490# 0.217f
C1377 a_n1500_45753# w_n1594_44514# 0.0172f
C1378 w_n1594_n28410# a_1500_n27074# 0.0023f
C1379 w_n1594_24738# a_n1500_23505# 0.0172f
C1380 a_n1500_n16047# a_n1500_n14811# 3.11f
C1381 a_1500_n45614# w_n1594_n44478# 0.0023f
C1382 a_n1558_23602# a_n1558_22366# 0.0105f
C1383 a_n1500_16089# a_1500_16186# 0.217f
C1384 w_n1594_n16050# a_n1558_n15950# 0.0187f
C1385 a_1500_42142# w_n1594_43278# 0.0023f
C1386 w_n1594_28446# a_n1558_27310# 0.0023f
C1387 a_n1500_n24699# a_n1558_n24602# 0.217f
C1388 w_n1594_n22230# a_n1500_n22227# 1.65f
C1389 a_1500_n23366# a_1500_n24602# 0.0105f
C1390 w_n1594_n60546# a_n1558_n60446# 0.0187f
C1391 a_1500_n61682# VSUBS 0.638f
C1392 a_n1558_n61682# VSUBS 0.638f
C1393 a_n1500_n61779# VSUBS 5.03f
C1394 a_1500_n60446# VSUBS 0.625f
C1395 a_n1558_n60446# VSUBS 0.625f
C1396 a_n1500_n60543# VSUBS 3.31f
C1397 a_1500_n59210# VSUBS 0.625f
C1398 a_n1558_n59210# VSUBS 0.625f
C1399 a_n1500_n59307# VSUBS 3.31f
C1400 a_1500_n57974# VSUBS 0.625f
C1401 a_n1558_n57974# VSUBS 0.625f
C1402 a_n1500_n58071# VSUBS 3.31f
C1403 a_1500_n56738# VSUBS 0.625f
C1404 a_n1558_n56738# VSUBS 0.625f
C1405 a_n1500_n56835# VSUBS 3.31f
C1406 a_1500_n55502# VSUBS 0.625f
C1407 a_n1558_n55502# VSUBS 0.625f
C1408 a_n1500_n55599# VSUBS 3.31f
C1409 a_1500_n54266# VSUBS 0.625f
C1410 a_n1558_n54266# VSUBS 0.625f
C1411 a_n1500_n54363# VSUBS 3.31f
C1412 a_1500_n53030# VSUBS 0.625f
C1413 a_n1558_n53030# VSUBS 0.625f
C1414 a_n1500_n53127# VSUBS 3.31f
C1415 a_1500_n51794# VSUBS 0.625f
C1416 a_n1558_n51794# VSUBS 0.625f
C1417 a_n1500_n51891# VSUBS 3.31f
C1418 a_1500_n50558# VSUBS 0.625f
C1419 a_n1558_n50558# VSUBS 0.625f
C1420 a_n1500_n50655# VSUBS 3.31f
C1421 a_1500_n49322# VSUBS 0.625f
C1422 a_n1558_n49322# VSUBS 0.625f
C1423 a_n1500_n49419# VSUBS 3.31f
C1424 a_1500_n48086# VSUBS 0.625f
C1425 a_n1558_n48086# VSUBS 0.625f
C1426 a_n1500_n48183# VSUBS 3.31f
C1427 a_1500_n46850# VSUBS 0.625f
C1428 a_n1558_n46850# VSUBS 0.625f
C1429 a_n1500_n46947# VSUBS 3.31f
C1430 a_1500_n45614# VSUBS 0.625f
C1431 a_n1558_n45614# VSUBS 0.625f
C1432 a_n1500_n45711# VSUBS 3.31f
C1433 a_1500_n44378# VSUBS 0.625f
C1434 a_n1558_n44378# VSUBS 0.625f
C1435 a_n1500_n44475# VSUBS 3.31f
C1436 a_1500_n43142# VSUBS 0.625f
C1437 a_n1558_n43142# VSUBS 0.625f
C1438 a_n1500_n43239# VSUBS 3.31f
C1439 a_1500_n41906# VSUBS 0.625f
C1440 a_n1558_n41906# VSUBS 0.625f
C1441 a_n1500_n42003# VSUBS 3.31f
C1442 a_1500_n40670# VSUBS 0.625f
C1443 a_n1558_n40670# VSUBS 0.625f
C1444 a_n1500_n40767# VSUBS 3.31f
C1445 a_1500_n39434# VSUBS 0.625f
C1446 a_n1558_n39434# VSUBS 0.625f
C1447 a_n1500_n39531# VSUBS 3.31f
C1448 a_1500_n38198# VSUBS 0.625f
C1449 a_n1558_n38198# VSUBS 0.625f
C1450 a_n1500_n38295# VSUBS 3.31f
C1451 a_1500_n36962# VSUBS 0.625f
C1452 a_n1558_n36962# VSUBS 0.625f
C1453 a_n1500_n37059# VSUBS 3.31f
C1454 a_1500_n35726# VSUBS 0.625f
C1455 a_n1558_n35726# VSUBS 0.625f
C1456 a_n1500_n35823# VSUBS 3.31f
C1457 a_1500_n34490# VSUBS 0.625f
C1458 a_n1558_n34490# VSUBS 0.625f
C1459 a_n1500_n34587# VSUBS 3.31f
C1460 a_1500_n33254# VSUBS 0.625f
C1461 a_n1558_n33254# VSUBS 0.625f
C1462 a_n1500_n33351# VSUBS 3.31f
C1463 a_1500_n32018# VSUBS 0.625f
C1464 a_n1558_n32018# VSUBS 0.625f
C1465 a_n1500_n32115# VSUBS 3.31f
C1466 a_1500_n30782# VSUBS 0.625f
C1467 a_n1558_n30782# VSUBS 0.625f
C1468 a_n1500_n30879# VSUBS 3.31f
C1469 a_1500_n29546# VSUBS 0.625f
C1470 a_n1558_n29546# VSUBS 0.625f
C1471 a_n1500_n29643# VSUBS 3.31f
C1472 a_1500_n28310# VSUBS 0.625f
C1473 a_n1558_n28310# VSUBS 0.625f
C1474 a_n1500_n28407# VSUBS 3.31f
C1475 a_1500_n27074# VSUBS 0.625f
C1476 a_n1558_n27074# VSUBS 0.625f
C1477 a_n1500_n27171# VSUBS 3.31f
C1478 a_1500_n25838# VSUBS 0.625f
C1479 a_n1558_n25838# VSUBS 0.625f
C1480 a_n1500_n25935# VSUBS 3.31f
C1481 a_1500_n24602# VSUBS 0.625f
C1482 a_n1558_n24602# VSUBS 0.625f
C1483 a_n1500_n24699# VSUBS 3.31f
C1484 a_1500_n23366# VSUBS 0.625f
C1485 a_n1558_n23366# VSUBS 0.625f
C1486 a_n1500_n23463# VSUBS 3.31f
C1487 a_1500_n22130# VSUBS 0.625f
C1488 a_n1558_n22130# VSUBS 0.625f
C1489 a_n1500_n22227# VSUBS 3.31f
C1490 a_1500_n20894# VSUBS 0.625f
C1491 a_n1558_n20894# VSUBS 0.625f
C1492 a_n1500_n20991# VSUBS 3.31f
C1493 a_1500_n19658# VSUBS 0.625f
C1494 a_n1558_n19658# VSUBS 0.625f
C1495 a_n1500_n19755# VSUBS 3.31f
C1496 a_1500_n18422# VSUBS 0.625f
C1497 a_n1558_n18422# VSUBS 0.625f
C1498 a_n1500_n18519# VSUBS 3.31f
C1499 a_1500_n17186# VSUBS 0.625f
C1500 a_n1558_n17186# VSUBS 0.625f
C1501 a_n1500_n17283# VSUBS 3.31f
C1502 a_1500_n15950# VSUBS 0.625f
C1503 a_n1558_n15950# VSUBS 0.625f
C1504 a_n1500_n16047# VSUBS 3.31f
C1505 a_1500_n14714# VSUBS 0.625f
C1506 a_n1558_n14714# VSUBS 0.625f
C1507 a_n1500_n14811# VSUBS 3.31f
C1508 a_1500_n13478# VSUBS 0.625f
C1509 a_n1558_n13478# VSUBS 0.625f
C1510 a_n1500_n13575# VSUBS 3.31f
C1511 a_1500_n12242# VSUBS 0.625f
C1512 a_n1558_n12242# VSUBS 0.625f
C1513 a_n1500_n12339# VSUBS 3.31f
C1514 a_1500_n11006# VSUBS 0.625f
C1515 a_n1558_n11006# VSUBS 0.625f
C1516 a_n1500_n11103# VSUBS 3.31f
C1517 a_1500_n9770# VSUBS 0.625f
C1518 a_n1558_n9770# VSUBS 0.625f
C1519 a_n1500_n9867# VSUBS 3.31f
C1520 a_1500_n8534# VSUBS 0.625f
C1521 a_n1558_n8534# VSUBS 0.625f
C1522 a_n1500_n8631# VSUBS 3.31f
C1523 a_1500_n7298# VSUBS 0.625f
C1524 a_n1558_n7298# VSUBS 0.625f
C1525 a_n1500_n7395# VSUBS 3.31f
C1526 a_1500_n6062# VSUBS 0.625f
C1527 a_n1558_n6062# VSUBS 0.625f
C1528 a_n1500_n6159# VSUBS 3.31f
C1529 a_1500_n4826# VSUBS 0.625f
C1530 a_n1558_n4826# VSUBS 0.625f
C1531 a_n1500_n4923# VSUBS 3.31f
C1532 a_1500_n3590# VSUBS 0.625f
C1533 a_n1558_n3590# VSUBS 0.625f
C1534 a_n1500_n3687# VSUBS 3.31f
C1535 a_1500_n2354# VSUBS 0.625f
C1536 a_n1558_n2354# VSUBS 0.625f
C1537 a_n1500_n2451# VSUBS 3.31f
C1538 a_1500_n1118# VSUBS 0.625f
C1539 a_n1558_n1118# VSUBS 0.625f
C1540 a_n1500_n1215# VSUBS 3.31f
C1541 a_1500_118# VSUBS 0.625f
C1542 a_n1558_118# VSUBS 0.625f
C1543 a_n1500_21# VSUBS 3.31f
C1544 a_1500_1354# VSUBS 0.625f
C1545 a_n1558_1354# VSUBS 0.625f
C1546 a_n1500_1257# VSUBS 3.31f
C1547 a_1500_2590# VSUBS 0.625f
C1548 a_n1558_2590# VSUBS 0.625f
C1549 a_n1500_2493# VSUBS 3.31f
C1550 a_1500_3826# VSUBS 0.625f
C1551 a_n1558_3826# VSUBS 0.625f
C1552 a_n1500_3729# VSUBS 3.31f
C1553 a_1500_5062# VSUBS 0.625f
C1554 a_n1558_5062# VSUBS 0.625f
C1555 a_n1500_4965# VSUBS 3.31f
C1556 a_1500_6298# VSUBS 0.625f
C1557 a_n1558_6298# VSUBS 0.625f
C1558 a_n1500_6201# VSUBS 3.31f
C1559 a_1500_7534# VSUBS 0.625f
C1560 a_n1558_7534# VSUBS 0.625f
C1561 a_n1500_7437# VSUBS 3.31f
C1562 a_1500_8770# VSUBS 0.625f
C1563 a_n1558_8770# VSUBS 0.625f
C1564 a_n1500_8673# VSUBS 3.31f
C1565 a_1500_10006# VSUBS 0.625f
C1566 a_n1558_10006# VSUBS 0.625f
C1567 a_n1500_9909# VSUBS 3.31f
C1568 a_1500_11242# VSUBS 0.625f
C1569 a_n1558_11242# VSUBS 0.625f
C1570 a_n1500_11145# VSUBS 3.31f
C1571 a_1500_12478# VSUBS 0.625f
C1572 a_n1558_12478# VSUBS 0.625f
C1573 a_n1500_12381# VSUBS 3.31f
C1574 a_1500_13714# VSUBS 0.625f
C1575 a_n1558_13714# VSUBS 0.625f
C1576 a_n1500_13617# VSUBS 3.31f
C1577 a_1500_14950# VSUBS 0.625f
C1578 a_n1558_14950# VSUBS 0.625f
C1579 a_n1500_14853# VSUBS 3.31f
C1580 a_1500_16186# VSUBS 0.625f
C1581 a_n1558_16186# VSUBS 0.625f
C1582 a_n1500_16089# VSUBS 3.31f
C1583 a_1500_17422# VSUBS 0.625f
C1584 a_n1558_17422# VSUBS 0.625f
C1585 a_n1500_17325# VSUBS 3.31f
C1586 a_1500_18658# VSUBS 0.625f
C1587 a_n1558_18658# VSUBS 0.625f
C1588 a_n1500_18561# VSUBS 3.31f
C1589 a_1500_19894# VSUBS 0.625f
C1590 a_n1558_19894# VSUBS 0.625f
C1591 a_n1500_19797# VSUBS 3.31f
C1592 a_1500_21130# VSUBS 0.625f
C1593 a_n1558_21130# VSUBS 0.625f
C1594 a_n1500_21033# VSUBS 3.31f
C1595 a_1500_22366# VSUBS 0.625f
C1596 a_n1558_22366# VSUBS 0.625f
C1597 a_n1500_22269# VSUBS 3.31f
C1598 a_1500_23602# VSUBS 0.625f
C1599 a_n1558_23602# VSUBS 0.625f
C1600 a_n1500_23505# VSUBS 3.31f
C1601 a_1500_24838# VSUBS 0.625f
C1602 a_n1558_24838# VSUBS 0.625f
C1603 a_n1500_24741# VSUBS 3.31f
C1604 a_1500_26074# VSUBS 0.625f
C1605 a_n1558_26074# VSUBS 0.625f
C1606 a_n1500_25977# VSUBS 3.31f
C1607 a_1500_27310# VSUBS 0.625f
C1608 a_n1558_27310# VSUBS 0.625f
C1609 a_n1500_27213# VSUBS 3.31f
C1610 a_1500_28546# VSUBS 0.625f
C1611 a_n1558_28546# VSUBS 0.625f
C1612 a_n1500_28449# VSUBS 3.31f
C1613 a_1500_29782# VSUBS 0.625f
C1614 a_n1558_29782# VSUBS 0.625f
C1615 a_n1500_29685# VSUBS 3.31f
C1616 a_1500_31018# VSUBS 0.625f
C1617 a_n1558_31018# VSUBS 0.625f
C1618 a_n1500_30921# VSUBS 3.31f
C1619 a_1500_32254# VSUBS 0.625f
C1620 a_n1558_32254# VSUBS 0.625f
C1621 a_n1500_32157# VSUBS 3.31f
C1622 a_1500_33490# VSUBS 0.625f
C1623 a_n1558_33490# VSUBS 0.625f
C1624 a_n1500_33393# VSUBS 3.31f
C1625 a_1500_34726# VSUBS 0.625f
C1626 a_n1558_34726# VSUBS 0.625f
C1627 a_n1500_34629# VSUBS 3.31f
C1628 a_1500_35962# VSUBS 0.625f
C1629 a_n1558_35962# VSUBS 0.625f
C1630 a_n1500_35865# VSUBS 3.31f
C1631 a_1500_37198# VSUBS 0.625f
C1632 a_n1558_37198# VSUBS 0.625f
C1633 a_n1500_37101# VSUBS 3.31f
C1634 a_1500_38434# VSUBS 0.625f
C1635 a_n1558_38434# VSUBS 0.625f
C1636 a_n1500_38337# VSUBS 3.31f
C1637 a_1500_39670# VSUBS 0.625f
C1638 a_n1558_39670# VSUBS 0.625f
C1639 a_n1500_39573# VSUBS 3.31f
C1640 a_1500_40906# VSUBS 0.625f
C1641 a_n1558_40906# VSUBS 0.625f
C1642 a_n1500_40809# VSUBS 3.31f
C1643 a_1500_42142# VSUBS 0.625f
C1644 a_n1558_42142# VSUBS 0.625f
C1645 a_n1500_42045# VSUBS 3.31f
C1646 a_1500_43378# VSUBS 0.625f
C1647 a_n1558_43378# VSUBS 0.625f
C1648 a_n1500_43281# VSUBS 3.31f
C1649 a_1500_44614# VSUBS 0.625f
C1650 a_n1558_44614# VSUBS 0.625f
C1651 a_n1500_44517# VSUBS 3.31f
C1652 a_1500_45850# VSUBS 0.625f
C1653 a_n1558_45850# VSUBS 0.625f
C1654 a_n1500_45753# VSUBS 3.31f
C1655 a_1500_47086# VSUBS 0.625f
C1656 a_n1558_47086# VSUBS 0.625f
C1657 a_n1500_46989# VSUBS 3.31f
C1658 a_1500_48322# VSUBS 0.625f
C1659 a_n1558_48322# VSUBS 0.625f
C1660 a_n1500_48225# VSUBS 3.31f
C1661 a_1500_49558# VSUBS 0.625f
C1662 a_n1558_49558# VSUBS 0.625f
C1663 a_n1500_49461# VSUBS 3.31f
C1664 a_1500_50794# VSUBS 0.625f
C1665 a_n1558_50794# VSUBS 0.625f
C1666 a_n1500_50697# VSUBS 3.31f
C1667 a_1500_52030# VSUBS 0.625f
C1668 a_n1558_52030# VSUBS 0.625f
C1669 a_n1500_51933# VSUBS 3.31f
C1670 a_1500_53266# VSUBS 0.625f
C1671 a_n1558_53266# VSUBS 0.625f
C1672 a_n1500_53169# VSUBS 3.31f
C1673 a_1500_54502# VSUBS 0.625f
C1674 a_n1558_54502# VSUBS 0.625f
C1675 a_n1500_54405# VSUBS 3.31f
C1676 a_1500_55738# VSUBS 0.625f
C1677 a_n1558_55738# VSUBS 0.625f
C1678 a_n1500_55641# VSUBS 3.31f
C1679 a_1500_56974# VSUBS 0.625f
C1680 a_n1558_56974# VSUBS 0.625f
C1681 a_n1500_56877# VSUBS 3.31f
C1682 a_1500_58210# VSUBS 0.625f
C1683 a_n1558_58210# VSUBS 0.625f
C1684 a_n1500_58113# VSUBS 3.31f
C1685 a_1500_59446# VSUBS 0.625f
C1686 a_n1558_59446# VSUBS 0.625f
C1687 a_n1500_59349# VSUBS 3.31f
C1688 a_1500_60682# VSUBS 0.638f
C1689 a_n1558_60682# VSUBS 0.638f
C1690 a_n1500_60585# VSUBS 5.03f
C1691 w_n1594_n61782# VSUBS 11.5f
C1692 w_n1594_n60546# VSUBS 11.5f
C1693 w_n1594_n59310# VSUBS 11.5f
C1694 w_n1594_n58074# VSUBS 11.5f
C1695 w_n1594_n56838# VSUBS 11.5f
C1696 w_n1594_n55602# VSUBS 11.5f
C1697 w_n1594_n54366# VSUBS 11.5f
C1698 w_n1594_n53130# VSUBS 11.5f
C1699 w_n1594_n51894# VSUBS 11.5f
C1700 w_n1594_n50658# VSUBS 11.5f
C1701 w_n1594_n49422# VSUBS 11.5f
C1702 w_n1594_n48186# VSUBS 11.5f
C1703 w_n1594_n46950# VSUBS 11.5f
C1704 w_n1594_n45714# VSUBS 11.5f
C1705 w_n1594_n44478# VSUBS 11.5f
C1706 w_n1594_n43242# VSUBS 11.5f
C1707 w_n1594_n42006# VSUBS 11.5f
C1708 w_n1594_n40770# VSUBS 11.5f
C1709 w_n1594_n39534# VSUBS 11.5f
C1710 w_n1594_n38298# VSUBS 11.5f
C1711 w_n1594_n37062# VSUBS 11.5f
C1712 w_n1594_n35826# VSUBS 11.5f
C1713 w_n1594_n34590# VSUBS 11.5f
C1714 w_n1594_n33354# VSUBS 11.5f
C1715 w_n1594_n32118# VSUBS 11.5f
C1716 w_n1594_n30882# VSUBS 11.5f
C1717 w_n1594_n29646# VSUBS 11.5f
C1718 w_n1594_n28410# VSUBS 11.5f
C1719 w_n1594_n27174# VSUBS 11.5f
C1720 w_n1594_n25938# VSUBS 11.5f
C1721 w_n1594_n24702# VSUBS 11.5f
C1722 w_n1594_n23466# VSUBS 11.5f
C1723 w_n1594_n22230# VSUBS 11.5f
C1724 w_n1594_n20994# VSUBS 11.5f
C1725 w_n1594_n19758# VSUBS 11.5f
C1726 w_n1594_n18522# VSUBS 11.5f
C1727 w_n1594_n17286# VSUBS 11.5f
C1728 w_n1594_n16050# VSUBS 11.5f
C1729 w_n1594_n14814# VSUBS 11.5f
C1730 w_n1594_n13578# VSUBS 11.5f
C1731 w_n1594_n12342# VSUBS 11.5f
C1732 w_n1594_n11106# VSUBS 11.5f
C1733 w_n1594_n9870# VSUBS 11.5f
C1734 w_n1594_n8634# VSUBS 11.5f
C1735 w_n1594_n7398# VSUBS 11.5f
C1736 w_n1594_n6162# VSUBS 11.5f
C1737 w_n1594_n4926# VSUBS 11.5f
C1738 w_n1594_n3690# VSUBS 11.5f
C1739 w_n1594_n2454# VSUBS 11.5f
C1740 w_n1594_n1218# VSUBS 11.5f
C1741 w_n1594_18# VSUBS 11.5f
C1742 w_n1594_1254# VSUBS 11.5f
C1743 w_n1594_2490# VSUBS 11.5f
C1744 w_n1594_3726# VSUBS 11.5f
C1745 w_n1594_4962# VSUBS 11.5f
C1746 w_n1594_6198# VSUBS 11.5f
C1747 w_n1594_7434# VSUBS 11.5f
C1748 w_n1594_8670# VSUBS 11.5f
C1749 w_n1594_9906# VSUBS 11.5f
C1750 w_n1594_11142# VSUBS 11.5f
C1751 w_n1594_12378# VSUBS 11.5f
C1752 w_n1594_13614# VSUBS 11.5f
C1753 w_n1594_14850# VSUBS 11.5f
C1754 w_n1594_16086# VSUBS 11.5f
C1755 w_n1594_17322# VSUBS 11.5f
C1756 w_n1594_18558# VSUBS 11.5f
C1757 w_n1594_19794# VSUBS 11.5f
C1758 w_n1594_21030# VSUBS 11.5f
C1759 w_n1594_22266# VSUBS 11.5f
C1760 w_n1594_23502# VSUBS 11.5f
C1761 w_n1594_24738# VSUBS 11.5f
C1762 w_n1594_25974# VSUBS 11.5f
C1763 w_n1594_27210# VSUBS 11.5f
C1764 w_n1594_28446# VSUBS 11.5f
C1765 w_n1594_29682# VSUBS 11.5f
C1766 w_n1594_30918# VSUBS 11.5f
C1767 w_n1594_32154# VSUBS 11.5f
C1768 w_n1594_33390# VSUBS 11.5f
C1769 w_n1594_34626# VSUBS 11.5f
C1770 w_n1594_35862# VSUBS 11.5f
C1771 w_n1594_37098# VSUBS 11.5f
C1772 w_n1594_38334# VSUBS 11.5f
C1773 w_n1594_39570# VSUBS 11.5f
C1774 w_n1594_40806# VSUBS 11.5f
C1775 w_n1594_42042# VSUBS 11.5f
C1776 w_n1594_43278# VSUBS 11.5f
C1777 w_n1594_44514# VSUBS 11.5f
C1778 w_n1594_45750# VSUBS 11.5f
C1779 w_n1594_46986# VSUBS 11.5f
C1780 w_n1594_48222# VSUBS 11.5f
C1781 w_n1594_49458# VSUBS 11.5f
C1782 w_n1594_50694# VSUBS 11.5f
C1783 w_n1594_51930# VSUBS 11.5f
C1784 w_n1594_53166# VSUBS 11.5f
C1785 w_n1594_54402# VSUBS 11.5f
C1786 w_n1594_55638# VSUBS 11.5f
C1787 w_n1594_56874# VSUBS 11.5f
C1788 w_n1594_58110# VSUBS 11.5f
C1789 w_n1594_59346# VSUBS 11.5f
C1790 w_n1594_60582# VSUBS 11.5f
.ends

.subckt sky130_fd_pr__nfet_01v8_WK8VRD a_n500_9156# a_n558_n10244# a_500_n2936# a_500_n5372#
+ a_n500_n1806# a_500_718# a_n500_3066# a_n500_n4242# a_n500_630# a_n500_n6678# a_n558_1936#
+ a_n558_4372# a_n558_n9026# a_n558_n6590# a_500_n500# a_500_6808# a_n500_6720# a_500_9244#
+ a_500_3154# a_500_n7808# a_n500_n9114# a_500_n4154# a_500_n1718# a_n558_n500# a_n500_n3024#
+ a_n558_6808# a_n558_9244# a_n558_n2936# a_n558_3154# a_n500_n10332# a_n558_n5372#
+ a_n558_718# a_n500_n588# a_n500_5502# a_500_8026# a_500_5590# a_n500_7938# a_500_n9026#
+ a_n500_1848# a_500_n6590# a_n500_4284# a_n500_n5460# a_n558_n7808# a_n500_n7896#
+ a_n558_8026# a_n558_n1718# a_n558_5590# a_n558_n4154# a_500_n10244# a_500_1936#
+ a_500_4372# VSUBS
X0 a_500_n10244# a_n500_n10332# a_n558_n10244# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X1 a_500_4372# a_n500_4284# a_n558_4372# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X2 a_500_n6590# a_n500_n6678# a_n558_n6590# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X3 a_500_5590# a_n500_5502# a_n558_5590# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X4 a_500_n1718# a_n500_n1806# a_n558_n1718# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X5 a_500_n2936# a_n500_n3024# a_n558_n2936# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X6 a_500_n4154# a_n500_n4242# a_n558_n4154# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X7 a_500_718# a_n500_630# a_n558_718# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X8 a_500_n5372# a_n500_n5460# a_n558_n5372# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X9 a_500_6808# a_n500_6720# a_n558_6808# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X10 a_500_8026# a_n500_7938# a_n558_8026# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X11 a_500_n500# a_n500_n588# a_n558_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X12 a_500_9244# a_n500_9156# a_n558_9244# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X13 a_500_1936# a_n500_1848# a_n558_1936# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X14 a_500_n7808# a_n500_n7896# a_n558_n7808# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X15 a_500_3154# a_n500_3066# a_n558_3154# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X16 a_500_n9026# a_n500_n9114# a_n558_n9026# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
C0 a_n558_718# a_n500_630# 0.204f
C1 a_n500_n4242# a_n500_n3024# 1.03f
C2 a_n500_n7896# a_n500_n6678# 1.03f
C3 a_n500_1848# a_n500_630# 1.03f
C4 a_n558_1936# a_500_1936# 0.0663f
C5 a_n558_3154# a_500_3154# 0.0663f
C6 a_500_4372# a_500_5590# 0.0113f
C7 a_n500_n588# a_n558_n500# 0.204f
C8 a_n500_4284# a_n558_4372# 0.204f
C9 a_n500_7938# a_500_8026# 0.204f
C10 a_n500_n588# a_n500_630# 1.03f
C11 a_n558_n10244# a_500_n10244# 0.0663f
C12 a_500_4372# a_n500_4284# 0.204f
C13 a_500_n5372# a_n500_n5460# 0.204f
C14 a_n500_n1806# a_500_n1718# 0.204f
C15 a_n500_n9114# a_n558_n9026# 0.204f
C16 a_n500_3066# a_n558_3154# 0.204f
C17 a_n558_3154# a_n558_1936# 0.0113f
C18 a_n500_n588# a_500_n500# 0.204f
C19 a_n500_n5460# a_n500_n6678# 1.03f
C20 a_n558_n1718# a_500_n1718# 0.0663f
C21 a_n500_5502# a_500_5590# 0.204f
C22 a_n558_n6590# a_n500_n6678# 0.204f
C23 a_500_n2936# a_500_n4154# 0.0113f
C24 a_n500_n4242# a_n558_n4154# 0.204f
C25 a_500_n9026# a_500_n10244# 0.0113f
C26 a_n558_n500# a_n558_n1718# 0.0113f
C27 a_n500_5502# a_n500_4284# 1.03f
C28 a_n500_6720# a_n500_7938# 1.03f
C29 a_n500_9156# a_n558_9244# 0.204f
C30 a_n500_n7896# a_n558_n7808# 0.204f
C31 a_n500_3066# a_500_3154# 0.204f
C32 a_n500_n4242# a_n500_n5460# 1.03f
C33 a_n558_n10244# a_n558_n9026# 0.0113f
C34 a_n500_5502# a_n500_6720# 1.03f
C35 a_n558_5590# a_n558_4372# 0.0113f
C36 a_n500_9156# a_n500_7938# 1.03f
C37 a_n558_9244# a_500_9244# 0.0663f
C38 a_n558_n2936# a_n500_n3024# 0.204f
C39 a_n558_n4154# a_500_n4154# 0.0663f
C40 a_n558_9244# a_n558_8026# 0.0113f
C41 a_n558_n7808# a_500_n7808# 0.0663f
C42 a_500_n2936# a_n500_n3024# 0.204f
C43 a_500_n7808# a_500_n9026# 0.0113f
C44 a_n500_3066# a_n500_4284# 1.03f
C45 a_n500_1848# a_500_1936# 0.204f
C46 a_n500_7938# a_n558_8026# 0.204f
C47 a_500_9244# a_500_8026# 0.0113f
C48 a_500_718# a_n500_630# 0.204f
C49 a_n558_n2936# a_500_n2936# 0.0663f
C50 a_n500_n10332# a_500_n10244# 0.204f
C51 a_n558_n7808# a_n558_n9026# 0.0113f
C52 a_n500_n9114# a_500_n9026# 0.204f
C53 a_500_n5372# a_500_n4154# 0.0113f
C54 a_500_n9026# a_n558_n9026# 0.0663f
C55 a_n558_n6590# a_n558_n7808# 0.0113f
C56 a_500_n500# a_500_n1718# 0.0113f
C57 a_500_6808# a_500_8026# 0.0113f
C58 a_n558_8026# a_500_8026# 0.0663f
C59 a_n500_n3024# a_n500_n1806# 1.03f
C60 a_500_718# a_500_n500# 0.0113f
C61 a_500_4372# a_n558_4372# 0.0663f
C62 a_500_n6590# a_500_n7808# 0.0113f
C63 a_n500_5502# a_n558_5590# 0.204f
C64 a_n558_n2936# a_n558_n4154# 0.0113f
C65 a_n558_n500# a_500_n500# 0.0663f
C66 a_500_6808# a_500_5590# 0.0113f
C67 a_n500_n588# a_n500_n1806# 1.03f
C68 a_n558_6808# a_n500_6720# 0.204f
C69 a_n558_3154# a_n558_4372# 0.0113f
C70 a_n558_n4154# a_n558_n5372# 0.0113f
C71 a_500_n5372# a_500_n6590# 0.0113f
C72 a_n558_n2936# a_n558_n1718# 0.0113f
C73 a_n558_n6590# a_500_n6590# 0.0663f
C74 a_n558_5590# a_500_5590# 0.0663f
C75 a_n500_n5460# a_n558_n5372# 0.204f
C76 a_n500_n9114# a_n500_n10332# 1.03f
C77 a_500_n6590# a_n500_n6678# 0.204f
C78 a_n500_n4242# a_500_n4154# 0.204f
C79 a_500_6808# a_n500_6720# 0.204f
C80 a_n500_9156# a_500_9244# 0.204f
C81 a_500_n5372# a_n558_n5372# 0.0663f
C82 a_n500_n7896# a_500_n7808# 0.204f
C83 a_n558_n5372# a_n558_n6590# 0.0113f
C84 a_500_3154# a_500_1936# 0.0113f
C85 a_n558_6808# a_500_6808# 0.0663f
C86 a_500_718# a_n558_718# 0.0663f
C87 a_n558_6808# a_n558_8026# 0.0113f
C88 a_n500_n7896# a_n500_n9114# 1.03f
C89 a_n500_3066# a_n500_1848# 1.03f
C90 a_n558_718# a_n558_1936# 0.0113f
C91 a_n500_1848# a_n558_1936# 0.204f
C92 a_500_3154# a_500_4372# 0.0113f
C93 a_500_n2936# a_500_n1718# 0.0113f
C94 a_n558_6808# a_n558_5590# 0.0113f
C95 a_n500_n1806# a_n558_n1718# 0.204f
C96 a_n558_n500# a_n558_718# 0.0113f
C97 a_500_718# a_500_1936# 0.0113f
C98 a_n500_n10332# a_n558_n10244# 0.204f
C99 a_500_n10244# VSUBS 0.581f
C100 a_n558_n10244# VSUBS 0.581f
C101 a_n500_n10332# VSUBS 2.28f
C102 a_500_n9026# VSUBS 0.571f
C103 a_n558_n9026# VSUBS 0.571f
C104 a_n500_n9114# VSUBS 1.71f
C105 a_500_n7808# VSUBS 0.571f
C106 a_n558_n7808# VSUBS 0.571f
C107 a_n500_n7896# VSUBS 1.71f
C108 a_500_n6590# VSUBS 0.571f
C109 a_n558_n6590# VSUBS 0.571f
C110 a_n500_n6678# VSUBS 1.71f
C111 a_500_n5372# VSUBS 0.571f
C112 a_n558_n5372# VSUBS 0.571f
C113 a_n500_n5460# VSUBS 1.71f
C114 a_500_n4154# VSUBS 0.571f
C115 a_n558_n4154# VSUBS 0.571f
C116 a_n500_n4242# VSUBS 1.71f
C117 a_500_n2936# VSUBS 0.571f
C118 a_n558_n2936# VSUBS 0.571f
C119 a_n500_n3024# VSUBS 1.71f
C120 a_500_n1718# VSUBS 0.571f
C121 a_n558_n1718# VSUBS 0.571f
C122 a_n500_n1806# VSUBS 1.71f
C123 a_500_n500# VSUBS 0.571f
C124 a_n558_n500# VSUBS 0.571f
C125 a_n500_n588# VSUBS 1.71f
C126 a_500_718# VSUBS 0.571f
C127 a_n558_718# VSUBS 0.571f
C128 a_n500_630# VSUBS 1.71f
C129 a_500_1936# VSUBS 0.571f
C130 a_n558_1936# VSUBS 0.571f
C131 a_n500_1848# VSUBS 1.71f
C132 a_500_3154# VSUBS 0.571f
C133 a_n558_3154# VSUBS 0.571f
C134 a_n500_3066# VSUBS 1.71f
C135 a_500_4372# VSUBS 0.571f
C136 a_n558_4372# VSUBS 0.571f
C137 a_n500_4284# VSUBS 1.71f
C138 a_500_5590# VSUBS 0.571f
C139 a_n558_5590# VSUBS 0.571f
C140 a_n500_5502# VSUBS 1.71f
C141 a_500_6808# VSUBS 0.571f
C142 a_n558_6808# VSUBS 0.571f
C143 a_n500_6720# VSUBS 1.71f
C144 a_500_8026# VSUBS 0.571f
C145 a_n558_8026# VSUBS 0.571f
C146 a_n500_7938# VSUBS 1.71f
C147 a_500_9244# VSUBS 0.581f
C148 a_n558_9244# VSUBS 0.581f
C149 a_n500_9156# VSUBS 2.28f
.ends

.subckt sky130_fd_pr__nfet_01v8_AH5E2K a_500_n500# a_n558_n500# a_n500_n588# VSUBS
X0 a_500_n500# a_n500_n588# a_n558_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
C0 a_n558_n500# a_500_n500# 0.0663f
C1 a_n500_n588# a_500_n500# 0.204f
C2 a_n500_n588# a_n558_n500# 0.204f
C3 a_500_n500# VSUBS 0.592f
C4 a_n558_n500# VSUBS 0.592f
C5 a_n500_n588# VSUBS 2.84f
.ends

.subckt sky130_fd_pr__pfet_01v8_C2U9V5 a_n300_n597# a_300_n500# w_n394_n600# a_n358_n500#
+ VSUBS
X0 a_300_n500# a_n300_n597# a_n358_n500# w_n394_n600# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=3
**devattr s=58000,2116 d=58000,2116
C0 a_n300_n597# a_n358_n500# 0.184f
C1 w_n394_n600# a_300_n500# 0.0187f
C2 a_n358_n500# a_300_n500# 0.107f
C3 w_n394_n600# a_n358_n500# 0.0187f
C4 a_n300_n597# a_300_n500# 0.184f
C5 w_n394_n600# a_n300_n597# 0.382f
C6 a_300_n500# VSUBS 0.548f
C7 a_n358_n500# VSUBS 0.548f
C8 a_n300_n597# VSUBS 1.42f
C9 w_n394_n600# VSUBS 2.84f
.ends

.subckt sky130_fd_pr__nfet_01v8_QP5WRD a_500_n2936# a_500_n5372# a_n500_n1806# a_500_718#
+ a_n500_3066# a_n500_n4242# a_n500_630# a_n500_n6678# a_n558_1936# a_n558_4372# a_n558_n9026#
+ a_n558_n6590# a_500_n500# a_500_6808# a_n500_6720# a_500_3154# a_500_n7808# a_n500_n9114#
+ a_500_n4154# a_500_n1718# a_n558_n500# a_n500_n3024# a_n558_6808# a_n558_n2936#
+ a_n558_3154# a_n558_n5372# a_n558_718# a_n500_n588# a_n500_5502# a_500_8026# a_500_5590#
+ a_n500_7938# a_500_n9026# a_n500_1848# a_500_n6590# a_n500_4284# a_n500_n5460# a_n558_n7808#
+ a_n500_n7896# a_n558_8026# a_n558_n1718# a_n558_5590# a_n558_n4154# a_500_1936#
+ a_500_4372# VSUBS
X0 a_500_4372# a_n500_4284# a_n558_4372# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X1 a_500_n6590# a_n500_n6678# a_n558_n6590# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X2 a_500_5590# a_n500_5502# a_n558_5590# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X3 a_500_n1718# a_n500_n1806# a_n558_n1718# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X4 a_500_n2936# a_n500_n3024# a_n558_n2936# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X5 a_500_n4154# a_n500_n4242# a_n558_n4154# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X6 a_500_718# a_n500_630# a_n558_718# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X7 a_500_n5372# a_n500_n5460# a_n558_n5372# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X8 a_500_6808# a_n500_6720# a_n558_6808# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X9 a_500_8026# a_n500_7938# a_n558_8026# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X10 a_500_n500# a_n500_n588# a_n558_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X11 a_500_1936# a_n500_1848# a_n558_1936# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X12 a_500_n7808# a_n500_n7896# a_n558_n7808# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X13 a_500_3154# a_n500_3066# a_n558_3154# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X14 a_500_n9026# a_n500_n9114# a_n558_n9026# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
C0 a_n558_n6590# a_n558_n7808# 0.0113f
C1 a_n500_6720# a_500_6808# 0.204f
C2 a_500_718# a_500_n500# 0.0113f
C3 a_n500_n7896# a_n500_n6678# 1.03f
C4 a_n500_n588# a_n558_n500# 0.204f
C5 a_n558_n2936# a_n558_n4154# 0.0113f
C6 a_500_3154# a_n500_3066# 0.204f
C7 a_n558_8026# a_500_8026# 0.0663f
C8 a_500_n500# a_500_n1718# 0.0113f
C9 a_n500_n1806# a_n558_n1718# 0.204f
C10 a_n500_n5460# a_500_n5372# 0.204f
C11 a_n500_4284# a_500_4372# 0.204f
C12 a_n558_718# a_500_718# 0.0663f
C13 a_n558_n500# a_n558_n1718# 0.0113f
C14 a_n558_n7808# a_500_n7808# 0.0663f
C15 a_n500_n1806# a_500_n1718# 0.204f
C16 a_n500_n4242# a_n558_n4154# 0.204f
C17 a_n558_n5372# a_500_n5372# 0.0663f
C18 a_n558_3154# a_n558_1936# 0.0113f
C19 a_n500_4284# a_n500_3066# 1.03f
C20 a_n500_7938# a_n500_6720# 1.03f
C21 a_n558_1936# a_n558_718# 0.0113f
C22 a_500_n5372# a_500_n6590# 0.0113f
C23 a_500_n2936# a_n558_n2936# 0.0663f
C24 a_n500_5502# a_n500_6720# 1.03f
C25 a_n558_4372# a_n558_3154# 0.0113f
C26 a_n500_4284# a_n500_5502# 1.03f
C27 a_n558_n6590# a_n500_n6678# 0.204f
C28 a_n558_8026# a_n558_6808# 0.0113f
C29 a_n500_n1806# a_n500_n3024# 1.03f
C30 a_n558_n6590# a_n558_n5372# 0.0113f
C31 a_500_1936# a_500_718# 0.0113f
C32 a_n500_630# a_n558_718# 0.204f
C33 a_n558_n5372# a_n558_n4154# 0.0113f
C34 a_n500_1848# a_500_1936# 0.204f
C35 a_500_8026# a_500_6808# 0.0113f
C36 a_n558_n1718# a_n558_n2936# 0.0113f
C37 a_n558_n6590# a_500_n6590# 0.0663f
C38 a_n500_n4242# a_n500_n5460# 1.03f
C39 a_n558_1936# a_500_1936# 0.0663f
C40 a_500_n5372# a_500_n4154# 0.0113f
C41 a_n500_6720# a_n558_6808# 0.204f
C42 a_n558_n9026# a_500_n9026# 0.0663f
C43 a_500_n7808# a_500_n6590# 0.0113f
C44 a_500_5590# a_500_6808# 0.0113f
C45 a_n500_4284# a_n558_4372# 0.204f
C46 a_n500_7938# a_500_8026# 0.204f
C47 a_n558_n500# a_500_n500# 0.0663f
C48 a_n500_n5460# a_n500_n6678# 1.03f
C49 a_n500_n5460# a_n558_n5372# 0.204f
C50 a_n558_6808# a_500_6808# 0.0663f
C51 a_500_n2936# a_500_n1718# 0.0113f
C52 a_n500_n3024# a_n558_n2936# 0.204f
C53 a_n500_3066# a_n500_1848# 1.03f
C54 a_500_3154# a_n558_3154# 0.0663f
C55 a_500_5590# a_500_4372# 0.0113f
C56 a_n558_n4154# a_500_n4154# 0.0663f
C57 a_n558_n500# a_n558_718# 0.0113f
C58 a_n558_5590# a_n500_5502# 0.204f
C59 a_n558_4372# a_500_4372# 0.0663f
C60 a_n558_n1718# a_500_n1718# 0.0663f
C61 a_n500_n4242# a_n500_n3024# 1.03f
C62 a_n500_n6678# a_500_n6590# 0.204f
C63 a_500_n2936# a_n500_n3024# 0.204f
C64 a_n500_n588# a_n500_630# 1.03f
C65 a_500_5590# a_n500_5502# 0.204f
C66 a_n558_n7808# a_n558_n9026# 0.0113f
C67 a_n500_n4242# a_500_n4154# 0.204f
C68 a_n500_n7896# a_n558_n7808# 0.204f
C69 a_500_n2936# a_500_n4154# 0.0113f
C70 a_n500_1848# a_n558_1936# 0.204f
C71 a_500_3154# a_500_1936# 0.0113f
C72 a_n558_5590# a_500_5590# 0.0663f
C73 a_n500_630# a_500_718# 0.204f
C74 a_n500_n7896# a_500_n7808# 0.204f
C75 a_n500_1848# a_n500_630# 1.03f
C76 a_n500_n9114# a_n558_n9026# 0.204f
C77 a_500_n7808# a_500_n9026# 0.0113f
C78 a_n558_5590# a_n558_6808# 0.0113f
C79 a_n500_n588# a_500_n500# 0.204f
C80 a_n558_5590# a_n558_4372# 0.0113f
C81 a_n500_n7896# a_n500_n9114# 1.03f
C82 a_n500_3066# a_n558_3154# 0.204f
C83 a_n500_n9114# a_500_n9026# 0.204f
C84 a_n500_n588# a_n500_n1806# 1.03f
C85 a_500_3154# a_500_4372# 0.0113f
C86 a_n500_7938# a_n558_8026# 0.204f
C87 a_500_n9026# VSUBS 0.581f
C88 a_n558_n9026# VSUBS 0.581f
C89 a_n500_n9114# VSUBS 2.28f
C90 a_500_n7808# VSUBS 0.571f
C91 a_n558_n7808# VSUBS 0.571f
C92 a_n500_n7896# VSUBS 1.71f
C93 a_500_n6590# VSUBS 0.571f
C94 a_n558_n6590# VSUBS 0.571f
C95 a_n500_n6678# VSUBS 1.71f
C96 a_500_n5372# VSUBS 0.571f
C97 a_n558_n5372# VSUBS 0.571f
C98 a_n500_n5460# VSUBS 1.71f
C99 a_500_n4154# VSUBS 0.571f
C100 a_n558_n4154# VSUBS 0.571f
C101 a_n500_n4242# VSUBS 1.71f
C102 a_500_n2936# VSUBS 0.571f
C103 a_n558_n2936# VSUBS 0.571f
C104 a_n500_n3024# VSUBS 1.71f
C105 a_500_n1718# VSUBS 0.571f
C106 a_n558_n1718# VSUBS 0.571f
C107 a_n500_n1806# VSUBS 1.71f
C108 a_500_n500# VSUBS 0.571f
C109 a_n558_n500# VSUBS 0.571f
C110 a_n500_n588# VSUBS 1.71f
C111 a_500_718# VSUBS 0.571f
C112 a_n558_718# VSUBS 0.571f
C113 a_n500_630# VSUBS 1.71f
C114 a_500_1936# VSUBS 0.571f
C115 a_n558_1936# VSUBS 0.571f
C116 a_n500_1848# VSUBS 1.71f
C117 a_500_3154# VSUBS 0.571f
C118 a_n558_3154# VSUBS 0.571f
C119 a_n500_3066# VSUBS 1.71f
C120 a_500_4372# VSUBS 0.571f
C121 a_n558_4372# VSUBS 0.571f
C122 a_n500_4284# VSUBS 1.71f
C123 a_500_5590# VSUBS 0.571f
C124 a_n558_5590# VSUBS 0.571f
C125 a_n500_5502# VSUBS 1.71f
C126 a_500_6808# VSUBS 0.571f
C127 a_n558_6808# VSUBS 0.571f
C128 a_n500_6720# VSUBS 1.71f
C129 a_500_8026# VSUBS 0.581f
C130 a_n558_8026# VSUBS 0.581f
C131 a_n500_7938# VSUBS 2.28f
.ends

.subckt sky130_fd_pr__pfet_01v8_UDM5A5 a_n558_n7916# a_n500_5583# a_500_1972# a_n558_8152#
+ a_n500_8055# a_500_4444# w_n594_3108# w_n594_6816# a_500_n2972# a_500_736# a_500_n5444#
+ a_n500_n597# w_n594_636# a_500_n500# w_n594_n3072# a_n558_1972# w_n594_n6780# w_n594_n600#
+ a_n500_1875# a_n558_4444# w_n594_n9252# a_n500_4347# a_n558_n6680# a_n558_n9152#
+ a_n500_n5541# a_n500_639# a_500_3208# a_n500_n8013# a_500_6916# a_500_n1736# a_n558_n500#
+ a_500_n4208# w_n594_5580# a_500_n7916# w_n594_8052# w_n594_n5544# a_n558_736# a_n558_3208#
+ w_n594_n8016# a_n558_n2972# a_n558_6916# a_n558_n5444# a_n500_n1833# a_n500_6819#
+ a_n500_n4305# w_n594_1872# a_500_5680# a_n500_n3069# w_n594_4344# a_n500_n6777#
+ a_500_8152# w_n594_n1836# a_n500_n9249# a_500_n6680# w_n594_n4308# a_n500_3111#
+ a_500_n9152# a_n558_n1736# a_n558_n4208# a_n558_5680# VSUBS
X0 a_500_1972# a_n500_1875# a_n558_1972# w_n594_1872# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X1 a_500_6916# a_n500_6819# a_n558_6916# w_n594_6816# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X2 a_500_4444# a_n500_4347# a_n558_4444# w_n594_4344# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X3 a_500_n9152# a_n500_n9249# a_n558_n9152# w_n594_n9252# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X4 a_500_3208# a_n500_3111# a_n558_3208# w_n594_3108# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X5 a_500_n2972# a_n500_n3069# a_n558_n2972# w_n594_n3072# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X6 a_500_n7916# a_n500_n8013# a_n558_n7916# w_n594_n8016# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X7 a_500_n5444# a_n500_n5541# a_n558_n5444# w_n594_n5544# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X8 a_500_n500# a_n500_n597# a_n558_n500# w_n594_n600# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X9 a_500_n1736# a_n500_n1833# a_n558_n1736# w_n594_n1836# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X10 a_500_n4208# a_n500_n4305# a_n558_n4208# w_n594_n4308# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X11 a_500_736# a_n500_639# a_n558_736# w_n594_636# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X12 a_500_n6680# a_n500_n6777# a_n558_n6680# w_n594_n6780# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X13 a_500_5680# a_n500_5583# a_n558_5680# w_n594_5580# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X14 a_500_8152# a_n500_8055# a_n558_8152# w_n594_8052# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
C0 w_n594_n600# a_n500_639# 0.00575f
C1 a_500_3208# w_n594_3108# 0.0187f
C2 a_n500_n4305# a_500_n4208# 0.204f
C3 w_n594_n6780# a_n500_n5541# 0.00575f
C4 a_n558_n7916# w_n594_n9252# 0.0023f
C5 a_500_n9152# w_n594_n9252# 0.0187f
C6 a_n500_n4305# w_n594_n3072# 0.00575f
C7 a_n558_n1736# a_n558_n500# 0.0105f
C8 a_500_736# w_n594_n600# 0.0023f
C9 w_n594_n9252# a_n500_n8013# 0.00575f
C10 w_n594_1872# a_n500_639# 0.00575f
C11 w_n594_n5544# a_500_n5444# 0.0187f
C12 a_n558_5680# w_n594_4344# 0.0023f
C13 a_n500_n5541# a_500_n5444# 0.204f
C14 a_n558_n1736# a_500_n1736# 0.0663f
C15 a_500_736# w_n594_1872# 0.0023f
C16 a_n500_4347# a_n500_3111# 1.03f
C17 a_n558_4444# a_500_4444# 0.0663f
C18 a_n500_n4305# w_n594_n4308# 0.593f
C19 a_500_5680# w_n594_4344# 0.0023f
C20 a_n558_736# w_n594_636# 0.0187f
C21 w_n594_n6780# a_500_n5444# 0.0023f
C22 a_500_8152# w_n594_8052# 0.0187f
C23 a_500_n6680# w_n594_n5544# 0.0023f
C24 a_n558_5680# a_n500_5583# 0.204f
C25 a_n558_3208# a_n558_1972# 0.0105f
C26 a_n558_n4208# a_n500_n4305# 0.204f
C27 a_n558_4444# a_n558_3208# 0.0105f
C28 a_n500_n1833# w_n594_n600# 0.00575f
C29 a_n558_736# a_n558_1972# 0.0105f
C30 a_n500_n597# w_n594_n600# 0.593f
C31 a_n558_4444# w_n594_5580# 0.0023f
C32 a_n500_1875# w_n594_1872# 0.593f
C33 a_n500_4347# w_n594_4344# 0.593f
C34 a_500_n7916# w_n594_n6780# 0.0023f
C35 a_500_5680# a_n500_5583# 0.204f
C36 a_n558_n2972# w_n594_n3072# 0.0187f
C37 a_500_8152# w_n594_6816# 0.0023f
C38 a_n558_6916# w_n594_8052# 0.0023f
C39 a_500_n6680# w_n594_n6780# 0.0187f
C40 w_n594_n5544# a_n558_n5444# 0.0187f
C41 a_500_736# a_500_n500# 0.0105f
C42 a_n500_n1833# w_n594_n1836# 0.593f
C43 a_n500_n597# w_n594_n1836# 0.00575f
C44 a_500_4444# w_n594_5580# 0.0023f
C45 a_n500_4347# w_n594_3108# 0.00575f
C46 a_n500_n5541# a_n558_n5444# 0.204f
C47 a_n500_n3069# w_n594_n3072# 0.593f
C48 a_n500_4347# a_n500_5583# 1.03f
C49 a_n558_n2972# w_n594_n4308# 0.0023f
C50 a_500_6916# w_n594_8052# 0.0023f
C51 a_n558_6916# w_n594_6816# 0.0187f
C52 a_500_n6680# a_500_n5444# 0.0105f
C53 w_n594_n5544# a_500_n4208# 0.0023f
C54 a_500_n9152# a_n500_n9249# 0.204f
C55 w_n594_1872# a_n558_1972# 0.0187f
C56 a_n500_n9249# a_n500_n8013# 1.03f
C57 w_n594_n6780# a_n558_n5444# 0.0023f
C58 a_500_4444# a_500_3208# 0.0105f
C59 a_500_n2972# w_n594_n1836# 0.0023f
C60 a_n500_3111# w_n594_4344# 0.00575f
C61 a_n500_n1833# a_n500_n3069# 1.03f
C62 a_n558_n4208# a_n558_n2972# 0.0105f
C63 a_n500_n3069# w_n594_n4308# 0.00575f
C64 a_500_n7916# a_500_n6680# 0.0105f
C65 a_n558_n2972# a_500_n2972# 0.0663f
C66 a_n558_n7916# a_n500_n8013# 0.204f
C67 a_n558_6916# w_n594_5580# 0.0023f
C68 a_500_6916# w_n594_6816# 0.0187f
C69 a_n558_n7916# a_n558_n6680# 0.0105f
C70 a_500_8152# a_500_6916# 0.0105f
C71 a_500_n1736# w_n594_n3072# 0.0023f
C72 w_n594_3108# a_500_1972# 0.0023f
C73 a_n558_3208# a_500_3208# 0.0663f
C74 a_n558_4444# a_n558_5680# 0.0105f
C75 a_n558_n5444# a_500_n5444# 0.0663f
C76 a_n558_n9152# w_n594_n9252# 0.0187f
C77 a_n500_n597# a_n558_n500# 0.204f
C78 a_n500_n597# a_500_n500# 0.204f
C79 a_500_736# a_500_1972# 0.0105f
C80 a_n500_3111# w_n594_3108# 0.593f
C81 a_n500_n3069# a_500_n2972# 0.204f
C82 a_n500_n9249# w_n594_n8016# 0.00575f
C83 a_n558_n500# w_n594_636# 0.0023f
C84 w_n594_636# a_500_n500# 0.0023f
C85 a_n500_8055# a_n558_8152# 0.204f
C86 w_n594_n4308# a_n500_n5541# 0.00575f
C87 a_500_6916# w_n594_5580# 0.0023f
C88 a_n558_n1736# w_n594_n3072# 0.0023f
C89 a_n558_736# w_n594_n600# 0.0023f
C90 a_n558_6916# a_500_6916# 0.0663f
C91 a_n500_6819# a_n500_5583# 1.03f
C92 a_n500_n8013# a_n500_n6777# 1.03f
C93 a_500_n4208# a_500_n5444# 0.0105f
C94 a_n558_n7916# w_n594_n8016# 0.0187f
C95 a_n500_n1833# a_500_n1736# 0.204f
C96 a_n558_n4208# w_n594_n5544# 0.0023f
C97 a_n500_n6777# a_n558_n6680# 0.204f
C98 a_500_n9152# w_n594_n8016# 0.0023f
C99 a_n558_5680# w_n594_6816# 0.0023f
C100 a_n558_3208# w_n594_1872# 0.0023f
C101 w_n594_n8016# a_n500_n8013# 0.593f
C102 w_n594_n8016# a_n558_n6680# 0.0023f
C103 a_n500_1875# a_500_1972# 0.204f
C104 a_n500_8055# a_n500_6819# 1.03f
C105 a_n558_736# w_n594_1872# 0.0023f
C106 a_n500_5583# w_n594_4344# 0.00575f
C107 a_n500_1875# a_n500_3111# 1.03f
C108 a_500_5680# a_500_4444# 0.0105f
C109 a_n500_4347# a_n558_4444# 0.204f
C110 a_n500_n1833# a_n558_n1736# 0.204f
C111 a_500_5680# w_n594_6816# 0.0023f
C112 a_500_n7916# w_n594_n9252# 0.0023f
C113 a_500_n1736# a_500_n2972# 0.0105f
C114 a_500_736# a_n500_639# 0.204f
C115 w_n594_n8016# a_n500_n6777# 0.00575f
C116 w_n594_n4308# a_500_n5444# 0.0023f
C117 a_500_3208# w_n594_1872# 0.0023f
C118 a_n558_5680# w_n594_5580# 0.0187f
C119 w_n594_636# a_500_1972# 0.0023f
C120 a_n558_5680# a_n558_6916# 0.0105f
C121 a_n500_4347# a_500_4444# 0.204f
C122 a_500_5680# w_n594_5580# 0.0187f
C123 a_n500_n3069# a_n500_n4305# 1.03f
C124 a_n558_1972# a_500_1972# 0.0663f
C125 a_n558_8152# w_n594_8052# 0.0187f
C126 a_n500_1875# a_n500_639# 1.03f
C127 a_n500_n4305# w_n594_n5544# 0.00575f
C128 a_n558_736# a_n558_n500# 0.0105f
C129 a_n500_1875# w_n594_3108# 0.00575f
C130 a_n500_4347# w_n594_5580# 0.00575f
C131 a_n558_n9152# a_n500_n9249# 0.204f
C132 a_n500_n4305# a_n500_n5541# 1.03f
C133 w_n594_n5544# a_n558_n6680# 0.0023f
C134 a_500_5680# a_500_6916# 0.0105f
C135 a_n558_n2972# w_n594_n1836# 0.0023f
C136 a_n500_n597# a_n500_639# 1.03f
C137 a_n500_6819# w_n594_8052# 0.00575f
C138 a_n558_8152# w_n594_6816# 0.0023f
C139 w_n594_636# a_n500_639# 0.593f
C140 a_n558_8152# a_500_8152# 0.0663f
C141 w_n594_n3072# a_500_n4208# 0.0023f
C142 a_n558_n7916# a_n558_n9152# 0.0105f
C143 a_n558_n7916# w_n594_n6780# 0.0023f
C144 w_n594_n4308# a_n558_n5444# 0.0023f
C145 a_n558_n9152# a_500_n9152# 0.0663f
C146 a_n558_n500# w_n594_n600# 0.0187f
C147 w_n594_n5544# a_n500_n6777# 0.00575f
C148 w_n594_n600# a_500_n500# 0.0187f
C149 w_n594_n6780# a_n500_n8013# 0.00575f
C150 a_n558_4444# w_n594_4344# 0.0187f
C151 a_n500_n3069# w_n594_n1836# 0.00575f
C152 a_500_736# w_n594_636# 0.0187f
C153 w_n594_n6780# a_n558_n6680# 0.0187f
C154 a_n500_n5541# a_n500_n6777# 1.03f
C155 a_n500_6819# w_n594_6816# 0.593f
C156 a_n500_n3069# a_n558_n2972# 0.204f
C157 a_n558_8152# a_n558_6916# 0.0105f
C158 a_n558_n4208# a_n558_n5444# 0.0105f
C159 w_n594_n4308# a_500_n4208# 0.0187f
C160 a_500_n1736# w_n594_n600# 0.0023f
C161 w_n594_3108# a_n558_1972# 0.0023f
C162 a_n500_3111# a_n558_3208# 0.204f
C163 a_500_5680# a_n558_5680# 0.0663f
C164 a_n500_n1833# w_n594_n3072# 0.00575f
C165 a_n558_n500# w_n594_n1836# 0.0023f
C166 w_n594_n1836# a_500_n500# 0.0023f
C167 w_n594_n6780# a_n500_n6777# 0.593f
C168 a_n558_4444# w_n594_3108# 0.0023f
C169 a_500_4444# w_n594_4344# 0.0187f
C170 a_n558_n9152# w_n594_n8016# 0.0023f
C171 a_n500_1875# w_n594_636# 0.00575f
C172 a_500_n7916# a_n558_n7916# 0.0663f
C173 a_n558_n4208# a_500_n4208# 0.0663f
C174 a_n500_6819# w_n594_5580# 0.00575f
C175 a_n558_n1736# w_n594_n600# 0.0023f
C176 a_500_n2972# a_500_n4208# 0.0105f
C177 a_500_n7916# a_500_n9152# 0.0105f
C178 a_500_3208# a_500_1972# 0.0105f
C179 a_n500_6819# a_n558_6916# 0.204f
C180 a_500_n7916# a_n500_n8013# 0.204f
C181 a_500_n1736# w_n594_n1836# 0.0187f
C182 a_n558_n4208# w_n594_n3072# 0.0023f
C183 a_n500_3111# a_500_3208# 0.204f
C184 a_500_n2972# w_n594_n3072# 0.0187f
C185 a_n500_n1833# a_n500_n597# 1.03f
C186 a_n558_3208# w_n594_4344# 0.0023f
C187 a_500_4444# w_n594_3108# 0.0023f
C188 a_n500_8055# w_n594_8052# 0.593f
C189 a_n500_n597# w_n594_636# 0.00575f
C190 a_n500_1875# a_n558_1972# 0.204f
C191 a_500_n6680# a_n558_n6680# 0.0663f
C192 a_n500_5583# w_n594_6816# 0.00575f
C193 a_n558_n1736# w_n594_n1836# 0.0187f
C194 a_n500_6819# a_500_6916# 0.204f
C195 a_n558_n4208# w_n594_n4308# 0.0187f
C196 w_n594_1872# a_500_1972# 0.0187f
C197 a_n558_n1736# a_n558_n2972# 0.0105f
C198 a_500_n2972# w_n594_n4308# 0.0023f
C199 a_n558_n500# a_500_n500# 0.0663f
C200 a_n558_736# a_n500_639# 0.204f
C201 a_n500_3111# w_n594_1872# 0.00575f
C202 a_500_3208# w_n594_4344# 0.0023f
C203 a_n558_3208# w_n594_3108# 0.0187f
C204 a_n500_8055# w_n594_6816# 0.00575f
C205 a_500_n7916# w_n594_n8016# 0.0187f
C206 w_n594_636# a_n558_1972# 0.0023f
C207 a_500_n6680# a_n500_n6777# 0.204f
C208 a_n500_8055# a_500_8152# 0.204f
C209 w_n594_n5544# a_n500_n5541# 0.593f
C210 a_n500_5583# w_n594_5580# 0.593f
C211 a_500_n6680# w_n594_n8016# 0.0023f
C212 a_n558_736# a_500_736# 0.0663f
C213 a_n558_n5444# a_n558_n6680# 0.0105f
C214 a_n500_n9249# w_n594_n9252# 0.593f
C215 a_500_n1736# a_500_n500# 0.0105f
C216 a_500_n9152# VSUBS 0.561f
C217 a_n558_n9152# VSUBS 0.561f
C218 a_n500_n9249# VSUBS 1.74f
C219 a_500_n7916# VSUBS 0.548f
C220 a_n558_n7916# VSUBS 0.548f
C221 a_n500_n8013# VSUBS 1.17f
C222 a_500_n6680# VSUBS 0.548f
C223 a_n558_n6680# VSUBS 0.548f
C224 a_n500_n6777# VSUBS 1.17f
C225 a_500_n5444# VSUBS 0.548f
C226 a_n558_n5444# VSUBS 0.548f
C227 a_n500_n5541# VSUBS 1.17f
C228 a_500_n4208# VSUBS 0.548f
C229 a_n558_n4208# VSUBS 0.548f
C230 a_n500_n4305# VSUBS 1.17f
C231 a_500_n2972# VSUBS 0.548f
C232 a_n558_n2972# VSUBS 0.548f
C233 a_n500_n3069# VSUBS 1.17f
C234 a_500_n1736# VSUBS 0.548f
C235 a_n558_n1736# VSUBS 0.548f
C236 a_n500_n1833# VSUBS 1.17f
C237 a_500_n500# VSUBS 0.548f
C238 a_n558_n500# VSUBS 0.548f
C239 a_n500_n597# VSUBS 1.17f
C240 a_500_736# VSUBS 0.548f
C241 a_n558_736# VSUBS 0.548f
C242 a_n500_639# VSUBS 1.17f
C243 a_500_1972# VSUBS 0.548f
C244 a_n558_1972# VSUBS 0.548f
C245 a_n500_1875# VSUBS 1.17f
C246 a_500_3208# VSUBS 0.548f
C247 a_n558_3208# VSUBS 0.548f
C248 a_n500_3111# VSUBS 1.17f
C249 a_500_4444# VSUBS 0.548f
C250 a_n558_4444# VSUBS 0.548f
C251 a_n500_4347# VSUBS 1.17f
C252 a_500_5680# VSUBS 0.548f
C253 a_n558_5680# VSUBS 0.548f
C254 a_n500_5583# VSUBS 1.17f
C255 a_500_6916# VSUBS 0.548f
C256 a_n558_6916# VSUBS 0.548f
C257 a_n500_6819# VSUBS 1.17f
C258 a_500_8152# VSUBS 0.561f
C259 a_n558_8152# VSUBS 0.561f
C260 a_n500_8055# VSUBS 1.74f
C261 w_n594_n9252# VSUBS 4.28f
C262 w_n594_n8016# VSUBS 4.28f
C263 w_n594_n6780# VSUBS 4.28f
C264 w_n594_n5544# VSUBS 4.28f
C265 w_n594_n4308# VSUBS 4.28f
C266 w_n594_n3072# VSUBS 4.28f
C267 w_n594_n1836# VSUBS 4.28f
C268 w_n594_n600# VSUBS 4.28f
C269 w_n594_636# VSUBS 4.28f
C270 w_n594_1872# VSUBS 4.28f
C271 w_n594_3108# VSUBS 4.28f
C272 w_n594_4344# VSUBS 4.28f
C273 w_n594_5580# VSUBS 4.28f
C274 w_n594_6816# VSUBS 4.28f
C275 w_n594_8052# VSUBS 4.28f
.ends

.subckt sky130_fd_pr__nfet_01v8_3ZAA45 a_100_n500# a_n158_n500# a_n100_n588# VSUBS
X0 a_100_n500# a_n100_n588# a_n158_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=1
**devattr s=58000,2116 d=58000,2116
C0 a_n100_n588# a_100_n500# 0.112f
C1 a_100_n500# a_n158_n500# 0.274f
C2 a_n100_n588# a_n158_n500# 0.112f
C3 a_100_n500# VSUBS 0.505f
C4 a_n158_n500# VSUBS 0.505f
C5 a_n100_n588# VSUBS 0.687f
.ends

.subckt sky130_fd_pr__pfet_01v8_SKU9VM a_n500_n597# a_500_n500# w_n594_n600# a_n558_n500#
+ VSUBS
X0 a_500_n500# a_n500_n597# a_n558_n500# w_n594_n600# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
C0 w_n594_n600# a_n558_n500# 0.0187f
C1 a_500_n500# a_n500_n597# 0.204f
C2 a_n558_n500# a_n500_n597# 0.204f
C3 a_n558_n500# a_500_n500# 0.0663f
C4 w_n594_n600# a_n500_n597# 0.593f
C5 w_n594_n600# a_500_n500# 0.0187f
C6 a_500_n500# VSUBS 0.573f
C7 a_n558_n500# VSUBS 0.573f
C8 a_n500_n597# VSUBS 2.31f
C9 w_n594_n600# VSUBS 4.28f
.ends

.subckt sky130_fd_pr__pfet_01v8_E769TZ a_n1558_11242# a_n1558_n14714# a_n1500_n43239#
+ w_n1594_n3690# a_n1500_n11103# a_n1558_50794# a_1500_n23366# a_n1500_n50655# w_n1594_n56838#
+ w_n1594_n24702# a_1500_n30782# a_n1500_3729# a_n1558_n60446# w_n1594_12378# w_n1594_n63018#
+ a_1500_n8534# a_n1558_14950# a_1500_n19658# a_n1500_n14811# a_n1500_n46947# w_n1594_9906#
+ w_n1594_n6162# a_1500_22366# a_n1500_22269# a_n1558_53266# a_n1558_n56738# a_n1558_n24602#
+ a_n1558_21130# a_n1500_n53127# w_n1594_n13578# a_n1558_60682# a_1500_n33254# a_n1500_n60543#
+ w_n1594_n20994# a_1500_n40670# a_1500_18658# a_n1558_49558# a_n1558_17422# w_n1594_22266#
+ a_n1500_n49419# w_n1594_n9870# a_n1500_25977# a_n1558_56974# a_n1500_n56835# a_1500_n29546#
+ a_n1558_n3590# a_1500_n36962# a_n1500_9909# a_n1558_n13478# a_1500_32254# a_n1500_32157#
+ a_n1558_n20894# a_n1500_n63015# w_n1594_18558# w_n1594_n23466# a_1500_n43142# w_n1594_n30882#
+ w_n1594_25974# a_n1500_n2451# a_1500_28546# a_1500_n7298# a_n1500_28449# a_n1558_59446#
+ a_n1558_27310# a_n1500_n13575# a_n1500_n59307# w_n1594_32154# w_n1594_n19758# a_1500_35962#
+ a_n1558_n6062# a_n1500_35865# a_1500_n39434# a_n1500_n20991# a_n1558_n23366# a_1500_n46850#
+ a_1500_42142# a_n1500_42045# a_n1558_n30782# w_n1594_n33354# w_n1594_28446# a_1500_n53030#
+ w_n1594_n40770# w_n1594_35862# a_n1558_n9770# w_n1594_18# a_n1558_16186# a_n1500_21#
+ a_n1558_n19658# a_n1500_n16047# a_1500_38434# a_n1500_38337# a_n1500_n55599# a_n1500_n23463#
+ w_n1594_n29646# a_1500_45850# w_n1594_42042# a_n1500_45753# a_n1558_40906# a_1500_n49322#
+ a_n1558_n33254# a_1500_52030# a_n1500_n8631# a_n1558_n40670# a_n1558_19894# w_n1594_n43242#
+ a_n1500_n19755# w_n1594_38334# w_n1594_45750# a_n1558_26074# a_n1558_n29546# a_1500_48322#
+ a_n1500_48225# a_1500_n38198# a_n1558_33490# a_n1558_n36962# a_n1500_n33351# w_n1594_n39534#
+ a_n1500_55641# a_1500_n59210# w_n1594_n46950# a_1500_n62918# a_n1558_n43142# a_n1558_29782#
+ w_n1594_n53130# a_n1500_n29643# w_n1594_48222# a_1500_37198# a_n1558_n39434# a_1500_58210#
+ a_n1500_58113# a_n1500_12381# a_1500_n1118# a_1500_n48086# a_n1558_n46850# a_1500_61918#
+ w_n1594_n49422# a_n1500_n7395# a_n1558_n53030# w_n1594_37098# a_n1558_39670# a_n1500_n39531#
+ w_n1594_58110# a_1500_n4826# w_n1594_61818# a_1500_47086# a_n1558_10006# a_n1558_n49322#
+ w_n1594_n2454# w_n1594_n38298# a_1500_2590# w_n1594_2490# w_n1594_n59310# a_n1500_6201#
+ a_n1500_18561# a_n1558_13714# a_n1558_2590# a_1500_n25838# a_n1558_n38198# a_1500_5062#
+ a_1500_118# a_n1558_n59210# w_n1594_n48186# w_n1594_n16050# a_n1558_n62918# a_1500_n32018#
+ a_n1500_2493# a_1500_24838# a_n1558_5062# a_n1500_n38295# w_n1594_n8634# a_1500_8770#
+ a_n1558_55738# a_n1558_23602# a_n1558_n2354# w_n1594_8670# a_1500_n35726# a_n1558_n48086#
+ a_1500_31018# w_n1594_n58074# w_n1594_24738# a_n1558_8770# a_n1500_n1215# a_n1558_12478#
+ a_n1500_n12339# a_n1500_n48183# a_1500_34726# a_n1500_34629# w_n1594_n25938# a_1500_n45614#
+ a_n1500_8673# w_n1594_n32118# a_n1500_n4923# w_n1594_34626# a_n1558_n8534# w_n1594_n7398#
+ a_n1558_22366# a_n1558_n25838# a_n1500_n22227# a_n1500_n58071# a_1500_44614# a_n1500_44517#
+ a_n1500_n61779# w_n1594_n35826# a_n1500_51933# a_1500_n55502# a_n1558_n32018# a_n1558_18658#
+ w_n1594_n42006# a_n1500_n18519# a_n1500_n25935# w_n1594_44514# w_n1594_51930# a_n1558_32254#
+ a_n1558_n35726# a_n1500_n32115# a_1500_54502# a_n1500_54405# a_1500_n44378# a_1500_n12242#
+ w_n1594_n45714# a_n1500_61821# a_1500_n51794# a_n1500_n3687# a_n1558_28546# a_n1558_n7298#
+ a_n1500_n28407# a_n1558_35962# a_n1500_n35823# w_n1594_54402# a_1500_n15950# a_1500_43378#
+ a_1500_11242# a_n1500_11145# a_n1558_42142# a_n1558_n45614# a_1500_50794# a_n1500_n42003#
+ a_n1500_50697# a_1500_n54266# a_1500_n22130# a_n1500_n6159# w_n1594_n55602# a_1500_n61682#
+ a_n1558_38434# a_n1500_n24699# w_n1594_43278# w_n1594_11142# a_1500_14950# a_n1500_46989#
+ a_n1558_45850# a_n1500_14853# a_1500_n18422# a_n1500_n45711# w_n1594_50694# a_1500_n57974#
+ a_n1500_n9867# w_n1594_n1218# a_1500_53266# a_1500_1354# a_n1500_53169# a_1500_21130#
+ a_n1500_21033# a_n1558_n55502# a_n1558_52030# w_n1594_1254# w_n1594_n12342# w_n1594_n44478#
+ a_1500_60682# a_n1500_60585# w_n1594_14850# w_n1594_n51894# w_n1594_46986# a_1500_49558#
+ a_1500_17422# a_n1558_48322# a_n1500_17325# a_n1500_n34587# a_1500_56974# a_n1558_1354#
+ w_n1594_53166# w_n1594_21030# w_n1594_n4926# a_n1500_56877# a_n1500_24741# a_1500_n3590#
+ a_1500_n28310# w_n1594_60582# w_n1594_4962# a_n1558_n44378# a_n1558_n12242# a_n1558_n51794#
+ w_n1594_17322# w_n1594_n22230# w_n1594_n54366# w_n1594_49458# a_n1500_1257# w_n1594_n61782#
+ w_n1594_56874# a_n1558_37198# a_n1500_n37059# a_1500_59446# a_1500_27310# a_1500_7534#
+ a_n1500_59349# a_n1500_27213# a_1500_n6062# a_1500_n17186# a_n1558_58210# a_n1558_n15950#
+ a_n1500_n44475# a_n1558_n1118# w_n1594_7434# w_n1594_n18522# a_n1558_61918# a_n1500_n51891#
+ a_n1558_n54266# a_1500_n41906# a_n1500_4965# a_n1558_n22130# a_n1558_n61682# w_n1594_59346#
+ w_n1594_27210# a_n1558_7534# a_1500_n9770# w_n1594_30918# a_n1558_n4826# a_1500_16186#
+ a_n1500_16089# a_n1558_47086# a_n1558_n18422# a_n1500_37101# a_n1558_n57974# a_1500_n27074#
+ a_n1500_n54363# a_1500_40906# w_n1594_n28410# a_n1500_40809# a_1500_n34490# a_n1500_7437#
+ w_n1594_16086# a_1500_19894# a_n1500_19797# w_n1594_40806# a_1500_26074# a_1500_6298#
+ a_n1558_n28310# w_n1594_6198# w_n1594_n17286# a_1500_33490# a_n1500_33393# w_n1594_19794#
+ a_n1558_6298# a_1500_29782# a_n1500_29685# a_n1558_24838# w_n1594_33390# a_n1558_n17186#
+ a_n1558_118# a_n1558_31018# w_n1594_n27174# a_n1500_43281# a_n1558_n41906# a_1500_n11006#
+ w_n1594_29682# w_n1594_n34590# a_1500_n50558# a_n1500_n17283# a_1500_39670# a_n1500_39573#
+ a_n1558_34726# a_1500_n14714# a_n1558_n27074# a_1500_10006# a_n1558_n34490# w_n1594_n37062#
+ w_n1594_39570# a_1500_n60446# a_n1500_n27171# a_1500_13714# a_n1500_13617# a_n1500_49461#
+ a_n1558_44614# a_n1500_n30879# a_1500_n56738# a_1500_n24602# w_n1594_n11106# w_n1594_n50658#
+ w_n1594_13614# a_1500_55738# a_1500_23602# a_1500_3826# a_n1500_23505# a_1500_n2354#
+ a_1500_n13478# a_n1558_54502# a_n1500_n40767# w_n1594_3726# w_n1594_n14814# a_n1500_30921#
+ a_1500_n20894# a_n1558_n11006# a_n1558_n50558# w_n1594_n60546# a_n1558_3826# w_n1594_55638#
+ w_n1594_23502# VSUBS a_1500_12478# a_n1558_43378#
X0 a_1500_53266# a_n1500_53169# a_n1558_53266# w_n1594_53166# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1 a_1500_n18422# a_n1500_n18519# a_n1558_n18422# w_n1594_n18522# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X2 a_1500_n45614# a_n1500_n45711# a_n1558_n45614# w_n1594_n45714# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X3 a_1500_n43142# a_n1500_n43239# a_n1558_n43142# w_n1594_n43242# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X4 a_1500_n22130# a_n1500_n22227# a_n1558_n22130# w_n1594_n22230# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X5 a_1500_n3590# a_n1500_n3687# a_n1558_n3590# w_n1594_n3690# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X6 a_1500_35962# a_n1500_35865# a_n1558_35962# w_n1594_35862# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X7 a_1500_33490# a_n1500_33393# a_n1558_33490# w_n1594_33390# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X8 a_1500_60682# a_n1500_60585# a_n1558_60682# w_n1594_60582# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X9 a_1500_12478# a_n1500_12381# a_n1558_12478# w_n1594_12378# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X10 a_1500_38434# a_n1500_38337# a_n1558_38434# w_n1594_38334# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X11 a_1500_6298# a_n1500_6201# a_n1558_6298# w_n1594_6198# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X12 a_1500_n55502# a_n1500_n55599# a_n1558_n55502# w_n1594_n55602# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X13 a_1500_n32018# a_n1500_n32115# a_n1558_n32018# w_n1594_n32118# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X14 a_1500_45850# a_n1500_45753# a_n1558_45850# w_n1594_45750# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X15 a_1500_24838# a_n1500_24741# a_n1558_24838# w_n1594_24738# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X16 a_1500_n38198# a_n1500_n38295# a_n1558_n38198# w_n1594_n38298# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X17 a_1500_22366# a_n1500_22269# a_n1558_22366# w_n1594_22266# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X18 a_1500_48322# a_n1500_48225# a_n1558_48322# w_n1594_48222# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X19 a_1500_n14714# a_n1500_n14811# a_n1558_n14714# w_n1594_n14814# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X20 a_1500_n41906# a_n1500_n42003# a_n1558_n41906# w_n1594_n42006# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X21 a_1500_n12242# a_n1500_n12339# a_n1558_n12242# w_n1594_n12342# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X22 a_1500_34726# a_n1500_34629# a_n1558_34726# w_n1594_34626# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X23 a_1500_61918# a_n1500_61821# a_n1558_61918# w_n1594_61818# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X24 a_1500_32254# a_n1500_32157# a_n1558_32254# w_n1594_32154# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X25 a_1500_n48086# a_n1500_n48183# a_n1558_n48086# w_n1594_n48186# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X26 a_1500_58210# a_n1500_58113# a_n1558_58210# w_n1594_58110# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X27 a_1500_n24602# a_n1500_n24699# a_n1558_n24602# w_n1594_n24702# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X28 a_1500_14950# a_n1500_14853# a_n1558_14950# w_n1594_14850# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X29 a_1500_n8534# a_n1500_n8631# a_n1558_n8534# w_n1594_n8634# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X30 a_1500_n57974# a_n1500_n58071# a_n1558_n57974# w_n1594_n58074# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X31 a_1500_n6062# a_n1500_n6159# a_n1558_n6062# w_n1594_n6162# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X32 a_1500_n34490# a_n1500_n34587# a_n1558_n34490# w_n1594_n34590# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X33 a_1500_17422# a_n1500_17325# a_n1558_17422# w_n1594_17322# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X34 a_1500_44614# a_n1500_44517# a_n1558_44614# w_n1594_44514# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X35 a_1500_42142# a_n1500_42045# a_n1558_42142# w_n1594_42042# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X36 a_1500_8770# a_n1500_8673# a_n1558_8770# w_n1594_8670# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X37 a_1500_n11006# a_n1500_n11103# a_n1558_n11006# w_n1594_n11106# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X38 a_1500_n19658# a_n1500_n19755# a_n1558_n19658# w_n1594_n19758# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X39 a_1500_n46850# a_n1500_n46947# a_n1558_n46850# w_n1594_n46950# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X40 a_1500_n17186# a_n1500_n17283# a_n1558_n17186# w_n1594_n17286# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X41 a_1500_27310# a_n1500_27213# a_n1558_27310# w_n1594_27210# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X42 a_1500_n44378# a_n1500_n44475# a_n1558_n44378# w_n1594_n44478# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X43 a_1500_54502# a_n1500_54405# a_n1558_54502# w_n1594_54402# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X44 a_1500_52030# a_n1500_51933# a_n1558_52030# w_n1594_51930# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X45 a_1500_31018# a_n1500_30921# a_n1558_31018# w_n1594_30918# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X46 a_1500_n4826# a_n1500_n4923# a_n1558_n4826# w_n1594_n4926# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X47 a_1500_37198# a_n1500_37101# a_n1558_37198# w_n1594_37098# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X48 a_1500_n2354# a_n1500_n2451# a_n1558_n2354# w_n1594_n2454# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X49 a_1500_n51794# a_n1500_n51891# a_n1558_n51794# w_n1594_n51894# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X50 a_1500_n29546# a_n1500_n29643# a_n1558_n29546# w_n1594_n29646# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X51 a_1500_13714# a_n1500_13617# a_n1558_13714# w_n1594_13614# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X52 a_1500_n56738# a_n1500_n56835# a_n1558_n56738# w_n1594_n56838# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X53 a_1500_11242# a_n1500_11145# a_n1558_11242# w_n1594_11142# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X54 a_1500_40906# a_n1500_40809# a_n1558_40906# w_n1594_40806# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X55 a_1500_n27074# a_n1500_n27171# a_n1558_n27074# w_n1594_n27174# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X56 a_1500_n54266# a_n1500_n54363# a_n1558_n54266# w_n1594_n54366# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X57 a_1500_19894# a_n1500_19797# a_n1558_19894# w_n1594_19794# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X58 a_1500_2590# a_n1500_2493# a_n1558_2590# w_n1594_2490# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X59 a_1500_n59210# a_n1500_n59307# a_n1558_n59210# w_n1594_n59310# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X60 a_1500_7534# a_n1500_7437# a_n1558_7534# w_n1594_7434# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X61 a_1500_49558# a_n1500_49461# a_n1558_49558# w_n1594_49458# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X62 a_1500_n36962# a_n1500_n37059# a_n1558_n36962# w_n1594_n37062# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X63 a_1500_5062# a_n1500_4965# a_n1558_5062# w_n1594_4962# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X64 a_1500_47086# a_n1500_46989# a_n1558_47086# w_n1594_46986# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X65 a_1500_n15950# a_n1500_n16047# a_n1558_n15950# w_n1594_n16050# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X66 a_1500_n61682# a_n1500_n61779# a_n1558_n61682# w_n1594_n61782# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X67 a_1500_n13478# a_n1500_n13575# a_n1558_n13478# w_n1594_n13578# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X68 a_1500_23602# a_n1500_23505# a_n1558_23602# w_n1594_23502# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X69 a_1500_n40670# a_n1500_n40767# a_n1558_n40670# w_n1594_n40770# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X70 a_1500_n39434# a_n1500_n39531# a_n1558_n39434# w_n1594_n39534# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X71 a_1500_21130# a_n1500_21033# a_n1558_21130# w_n1594_21030# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X72 a_1500_29782# a_n1500_29685# a_n1558_29782# w_n1594_29682# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X73 a_1500_56974# a_n1500_56877# a_n1558_56974# w_n1594_56874# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X74 a_1500_59446# a_n1500_59349# a_n1558_59446# w_n1594_59346# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X75 a_1500_n20894# a_n1500_n20991# a_n1558_n20894# w_n1594_n20994# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X76 a_1500_n25838# a_n1500_n25935# a_n1558_n25838# w_n1594_n25938# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X77 a_1500_n23366# a_n1500_n23463# a_n1558_n23366# w_n1594_n23466# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X78 a_1500_n50558# a_n1500_n50655# a_n1558_n50558# w_n1594_n50658# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X79 a_1500_n49322# a_n1500_n49419# a_n1558_n49322# w_n1594_n49422# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X80 a_1500_n1118# a_n1500_n1215# a_n1558_n1118# w_n1594_n1218# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X81 a_1500_n9770# a_n1500_n9867# a_n1558_n9770# w_n1594_n9870# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X82 a_1500_n28310# a_n1500_n28407# a_n1558_n28310# w_n1594_n28410# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X83 a_1500_n7298# a_n1500_n7395# a_n1558_n7298# w_n1594_n7398# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X84 a_1500_10006# a_n1500_9909# a_n1558_10006# w_n1594_9906# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X85 a_1500_39670# a_n1500_39573# a_n1558_39670# w_n1594_39570# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X86 a_1500_18658# a_n1500_18561# a_n1558_18658# w_n1594_18558# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X87 a_1500_n53030# a_n1500_n53127# a_n1558_n53030# w_n1594_n53130# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X88 a_1500_3826# a_n1500_3729# a_n1558_3826# w_n1594_3726# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X89 a_1500_16186# a_n1500_16089# a_n1558_16186# w_n1594_16086# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X90 a_1500_1354# a_n1500_1257# a_n1558_1354# w_n1594_1254# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X91 a_1500_43378# a_n1500_43281# a_n1558_43378# w_n1594_43278# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X92 a_1500_n30782# a_n1500_n30879# a_n1558_n30782# w_n1594_n30882# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X93 a_1500_118# a_n1500_21# a_n1558_118# w_n1594_18# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X94 a_1500_n35726# a_n1500_n35823# a_n1558_n35726# w_n1594_n35826# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X95 a_1500_n62918# a_n1500_n63015# a_n1558_n62918# w_n1594_n63018# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X96 a_1500_n33254# a_n1500_n33351# a_n1558_n33254# w_n1594_n33354# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X97 a_1500_n60446# a_n1500_n60543# a_n1558_n60446# w_n1594_n60546# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X98 a_1500_50794# a_n1500_50697# a_n1558_50794# w_n1594_50694# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X99 a_1500_28546# a_n1500_28449# a_n1558_28546# w_n1594_28446# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X100 a_1500_55738# a_n1500_55641# a_n1558_55738# w_n1594_55638# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X101 a_1500_26074# a_n1500_25977# a_n1558_26074# w_n1594_25974# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
C0 w_n1594_n30882# a_n1500_n29643# 0.0172f
C1 a_1500_n2354# w_n1594_n1218# 0.0023f
C2 a_n1500_n4923# w_n1594_n6162# 0.0172f
C3 a_1500_19894# a_n1500_19797# 0.217f
C4 a_n1558_33490# w_n1594_34626# 0.0023f
C5 a_n1500_39573# w_n1594_40806# 0.0172f
C6 a_n1500_25977# a_n1500_24741# 3.11f
C7 w_n1594_n55602# a_1500_n55502# 0.0187f
C8 a_n1500_n32115# a_n1500_n30879# 3.11f
C9 w_n1594_23502# a_n1500_22269# 0.0172f
C10 a_1500_42142# a_n1500_42045# 0.217f
C11 a_1500_18658# w_n1594_17322# 0.0023f
C12 w_n1594_4962# a_1500_5062# 0.0187f
C13 a_n1500_46989# a_n1500_48225# 3.11f
C14 a_n1500_n29643# w_n1594_n28410# 0.0172f
C15 a_1500_n6062# w_n1594_n7398# 0.0023f
C16 a_n1558_27310# w_n1594_28446# 0.0023f
C17 a_n1500_59349# a_n1500_58113# 3.11f
C18 a_n1558_n25838# a_n1558_n27074# 0.0105f
C19 a_n1558_21130# w_n1594_22266# 0.0023f
C20 a_1500_n54266# w_n1594_n53130# 0.0023f
C21 a_n1558_32254# w_n1594_30918# 0.0023f
C22 a_n1500_n16047# w_n1594_n16050# 1.65f
C23 a_1500_n3590# w_n1594_n3690# 0.0187f
C24 a_1500_n59210# a_1500_n57974# 0.0105f
C25 a_1500_12478# w_n1594_12378# 0.0187f
C26 a_n1500_38337# a_n1558_38434# 0.217f
C27 a_n1558_n36962# a_n1558_n38198# 0.0105f
C28 a_1500_26074# w_n1594_25974# 0.0187f
C29 a_1500_17422# w_n1594_16086# 0.0023f
C30 a_n1558_n45614# w_n1594_n45714# 0.0187f
C31 w_n1594_58110# a_n1500_59349# 0.0172f
C32 a_1500_n6062# w_n1594_n4926# 0.0023f
C33 a_n1500_13617# a_1500_13714# 0.217f
C34 a_1500_n41906# w_n1594_n40770# 0.0023f
C35 w_n1594_n61782# a_1500_n62918# 0.0023f
C36 a_n1558_38434# a_n1558_37198# 0.0105f
C37 a_n1558_n13478# w_n1594_n14814# 0.0023f
C38 a_n1500_17325# w_n1594_17322# 1.65f
C39 a_1500_n19658# w_n1594_n20994# 0.0023f
C40 a_n1500_35865# w_n1594_37098# 0.0172f
C41 w_n1594_n59310# a_1500_n57974# 0.0023f
C42 w_n1594_n18522# a_n1558_n18422# 0.0187f
C43 a_1500_n7298# w_n1594_n7398# 0.0187f
C44 w_n1594_55638# a_n1558_56974# 0.0023f
C45 a_1500_12478# a_n1500_12381# 0.217f
C46 a_n1558_n25838# w_n1594_n25938# 0.0187f
C47 a_1500_n23366# w_n1594_n24702# 0.0023f
C48 a_n1500_n45711# w_n1594_n44478# 0.0172f
C49 a_n1500_n6159# w_n1594_n6162# 1.65f
C50 a_n1558_n46850# w_n1594_n48186# 0.0023f
C51 w_n1594_n28410# a_1500_n27074# 0.0023f
C52 w_n1594_n27174# a_n1500_n28407# 0.0172f
C53 a_n1500_21# a_1500_118# 0.217f
C54 a_n1558_n4826# a_n1500_n4923# 0.217f
C55 a_1500_n17186# w_n1594_n16050# 0.0023f
C56 a_1500_27310# w_n1594_27210# 0.0187f
C57 a_n1558_7534# a_n1558_8770# 0.0105f
C58 a_n1558_29782# w_n1594_29682# 0.0187f
C59 a_n1500_n61779# a_1500_n61682# 0.217f
C60 a_n1558_32254# w_n1594_33390# 0.0023f
C61 w_n1594_n58074# a_1500_n59210# 0.0023f
C62 w_n1594_n30882# a_n1500_n32115# 0.0172f
C63 a_n1558_18658# w_n1594_18558# 0.0187f
C64 a_1500_56974# a_1500_58210# 0.0105f
C65 a_1500_n19658# w_n1594_n18522# 0.0023f
C66 w_n1594_n60546# a_1500_n61682# 0.0023f
C67 a_n1558_n13478# a_n1500_n13575# 0.217f
C68 a_n1558_27310# w_n1594_25974# 0.0023f
C69 a_1500_45850# w_n1594_45750# 0.0187f
C70 a_n1500_n32115# a_n1500_n33351# 3.11f
C71 a_1500_n28310# a_n1500_n28407# 0.217f
C72 w_n1594_9906# a_n1500_11145# 0.0172f
C73 w_n1594_56874# a_1500_56974# 0.0187f
C74 a_n1558_n48086# w_n1594_n49422# 0.0023f
C75 w_n1594_58110# a_1500_59446# 0.0023f
C76 a_1500_28546# w_n1594_27210# 0.0023f
C77 a_n1558_40906# a_n1558_39670# 0.0105f
C78 a_n1500_n55599# a_n1500_n56835# 3.11f
C79 a_n1500_21# a_n1500_1257# 3.11f
C80 a_n1558_56974# a_n1558_55738# 0.0105f
C81 a_1500_13714# a_1500_14950# 0.0105f
C82 a_1500_35962# w_n1594_34626# 0.0023f
C83 a_1500_48322# w_n1594_49458# 0.0023f
C84 a_1500_n41906# a_1500_n43142# 0.0105f
C85 a_n1500_n43239# a_n1558_n43142# 0.217f
C86 a_n1500_61821# a_n1558_61918# 0.217f
C87 a_n1558_50794# w_n1594_50694# 0.0187f
C88 w_n1594_54402# a_1500_54502# 0.0187f
C89 a_n1558_44614# a_n1558_45850# 0.0105f
C90 w_n1594_n55602# a_1500_n54266# 0.0023f
C91 a_1500_n3590# a_1500_n4826# 0.0105f
C92 w_n1594_3726# a_n1558_3826# 0.0187f
C93 a_n1500_n50655# w_n1594_n51894# 0.0172f
C94 a_1500_19894# w_n1594_18558# 0.0023f
C95 w_n1594_60582# a_n1558_61918# 0.0023f
C96 w_n1594_14850# a_n1558_14950# 0.0187f
C97 w_n1594_23502# a_n1500_24741# 0.0172f
C98 a_n1558_118# a_n1558_n1118# 0.0105f
C99 a_n1558_18658# w_n1594_19794# 0.0023f
C100 a_n1500_42045# a_n1500_40809# 3.11f
C101 a_n1558_n28310# w_n1594_n27174# 0.0023f
C102 a_n1500_7437# a_1500_7534# 0.217f
C103 a_n1500_n23463# w_n1594_n24702# 0.0172f
C104 a_n1558_1354# a_n1558_118# 0.0105f
C105 a_n1500_n25935# a_1500_n25838# 0.217f
C106 w_n1594_2490# a_n1500_1257# 0.0172f
C107 a_n1558_31018# w_n1594_32154# 0.0023f
C108 a_1500_2590# w_n1594_3726# 0.0023f
C109 a_n1500_32157# w_n1594_32154# 1.65f
C110 a_1500_n53030# w_n1594_n53130# 0.0187f
C111 a_n1558_n34490# w_n1594_n33354# 0.0023f
C112 a_1500_n14714# a_n1500_n14811# 0.217f
C113 w_n1594_6198# a_n1500_4965# 0.0172f
C114 a_n1500_n37059# a_1500_n36962# 0.217f
C115 a_n1558_n15950# w_n1594_n16050# 0.0187f
C116 a_n1558_n23366# a_n1558_n22130# 0.0105f
C117 w_n1594_n58074# a_n1500_n59307# 0.0172f
C118 w_n1594_n54366# a_n1500_n55599# 0.0172f
C119 a_1500_27310# w_n1594_28446# 0.0023f
C120 w_n1594_59346# a_n1500_60585# 0.0172f
C121 a_1500_39670# w_n1594_40806# 0.0023f
C122 w_n1594_n7398# a_n1500_n8631# 0.0172f
C123 a_n1558_n44378# w_n1594_n45714# 0.0023f
C124 w_n1594_n43242# a_1500_n43142# 0.0187f
C125 a_1500_49558# a_1500_50794# 0.0105f
C126 a_1500_n40670# w_n1594_n39534# 0.0023f
C127 a_1500_n40670# w_n1594_n40770# 0.0187f
C128 w_n1594_n61782# a_1500_n61682# 0.0187f
C129 a_1500_19894# w_n1594_19794# 0.0187f
C130 a_1500_n9770# w_n1594_n9870# 0.0187f
C131 w_n1594_n17286# a_n1558_n18422# 0.0023f
C132 a_n1558_n24602# w_n1594_n25938# 0.0023f
C133 a_n1558_8770# a_n1558_10006# 0.0105f
C134 w_n1594_28446# a_1500_28546# 0.0187f
C135 a_1500_n30782# w_n1594_n32118# 0.0023f
C136 a_n1500_38337# a_1500_38434# 0.217f
C137 a_1500_n7298# a_1500_n6062# 0.0105f
C138 a_n1500_55641# a_n1500_54405# 3.11f
C139 a_1500_n13478# w_n1594_n14814# 0.0023f
C140 a_1500_n48086# w_n1594_n46950# 0.0023f
C141 w_n1594_n27174# a_n1500_n27171# 1.65f
C142 a_n1500_n51891# a_n1558_n51794# 0.217f
C143 a_1500_21130# w_n1594_19794# 0.0023f
C144 w_n1594_2490# a_n1500_2493# 1.65f
C145 a_n1558_n60446# a_n1558_n61682# 0.0105f
C146 w_n1594_n60546# a_1500_n60446# 0.0187f
C147 a_1500_11242# w_n1594_9906# 0.0023f
C148 a_n1500_38337# w_n1594_39570# 0.0172f
C149 a_1500_n38198# w_n1594_n39534# 0.0023f
C150 a_1500_48322# a_1500_47086# 0.0105f
C151 a_1500_n22130# w_n1594_n22230# 0.0187f
C152 w_n1594_n63018# a_1500_n62918# 0.0187f
C153 a_n1500_n46947# a_n1558_n46850# 0.217f
C154 a_1500_38434# a_1500_37198# 0.0105f
C155 a_1500_n45614# a_1500_n46850# 0.0105f
C156 a_n1558_n28310# a_n1558_n27074# 0.0105f
C157 a_1500_n13478# a_n1500_n13575# 0.217f
C158 w_n1594_n50658# a_n1500_n51891# 0.0172f
C159 w_n1594_56874# a_n1500_56877# 1.65f
C160 a_n1558_38434# a_n1558_39670# 0.0105f
C161 a_n1500_24741# w_n1594_25974# 0.0172f
C162 a_1500_27310# w_n1594_25974# 0.0023f
C163 a_n1558_n17186# a_n1558_n15950# 0.0105f
C164 w_n1594_n34590# a_n1558_n34490# 0.0187f
C165 w_n1594_n11106# a_n1558_n9770# 0.0023f
C166 a_n1500_35865# a_1500_35962# 0.217f
C167 a_1500_n24602# w_n1594_n24702# 0.0187f
C168 a_n1500_9909# w_n1594_9906# 1.65f
C169 a_n1500_n9867# w_n1594_n8634# 0.0172f
C170 a_1500_50794# w_n1594_50694# 0.0187f
C171 a_n1500_35865# a_n1500_37101# 3.11f
C172 w_n1594_56874# a_n1500_55641# 0.0172f
C173 w_n1594_59346# a_n1558_59446# 0.0187f
C174 w_n1594_37098# a_1500_35962# 0.0023f
C175 w_n1594_48222# a_1500_47086# 0.0023f
C176 a_n1500_34629# w_n1594_34626# 1.65f
C177 a_n1558_50794# w_n1594_49458# 0.0023f
C178 a_1500_11242# a_1500_12478# 0.0105f
C179 a_n1500_n34587# w_n1594_n35826# 0.0172f
C180 a_1500_48322# w_n1594_46986# 0.0023f
C181 w_n1594_1254# a_1500_118# 0.0023f
C182 a_n1500_37101# w_n1594_37098# 1.65f
C183 w_n1594_2490# a_1500_1354# 0.0023f
C184 a_n1500_13617# w_n1594_12378# 0.0172f
C185 a_n1500_n38295# w_n1594_n37062# 0.0172f
C186 a_1500_8770# w_n1594_9906# 0.0023f
C187 w_n1594_54402# a_n1500_53169# 0.0172f
C188 w_n1594_n19758# a_1500_n18422# 0.0023f
C189 a_n1500_n7395# w_n1594_n8634# 0.0172f
C190 a_n1500_n24699# w_n1594_n23466# 0.0172f
C191 w_n1594_61818# a_1500_61918# 0.0187f
C192 a_n1500_51933# a_n1500_53169# 3.11f
C193 a_n1558_n33254# w_n1594_n33354# 0.0187f
C194 w_n1594_n56838# a_n1500_n58071# 0.0172f
C195 a_1500_n33254# w_n1594_n32118# 0.0023f
C196 a_1500_n25838# a_1500_n27074# 0.0105f
C197 a_1500_n51794# w_n1594_n53130# 0.0023f
C198 a_n1500_n27171# a_n1558_n27074# 0.217f
C199 a_n1558_43378# w_n1594_43278# 0.0187f
C200 w_n1594_58110# a_n1558_56974# 0.0023f
C201 a_n1558_n35726# a_n1558_n36962# 0.0105f
C202 w_n1594_n54366# a_n1500_n54363# 1.65f
C203 a_n1500_42045# a_n1558_42142# 0.217f
C204 a_n1500_12381# w_n1594_11142# 0.0172f
C205 a_1500_n44378# a_1500_n43142# 0.0105f
C206 a_n1558_n44378# a_n1500_n44475# 0.217f
C207 a_n1500_6201# a_n1500_4965# 3.11f
C208 a_n1558_13714# a_n1558_14950# 0.0105f
C209 a_n1500_n30879# w_n1594_n29646# 0.0172f
C210 w_n1594_n42006# a_n1500_n43239# 0.0172f
C211 w_n1594_n43242# a_1500_n41906# 0.0023f
C212 a_1500_n39434# w_n1594_n39534# 0.0187f
C213 a_n1558_n22130# a_n1558_n20894# 0.0105f
C214 a_1500_n39434# w_n1594_n40770# 0.0023f
C215 a_n1558_n11006# w_n1594_n9870# 0.0023f
C216 a_1500_22366# w_n1594_23502# 0.0023f
C217 a_n1500_n4923# w_n1594_n3690# 0.0172f
C218 w_n1594_1254# a_n1500_1257# 1.65f
C219 a_n1500_3729# a_n1500_4965# 3.11f
C220 a_n1500_13617# a_n1500_12381# 3.11f
C221 w_n1594_n61782# a_1500_n60446# 0.0023f
C222 a_n1500_49461# a_n1500_50697# 3.11f
C223 w_n1594_22266# a_n1500_22269# 1.65f
C224 w_n1594_n9870# a_n1500_n8631# 0.0172f
C225 a_1500_n46850# w_n1594_n46950# 0.0187f
C226 w_n1594_n25938# a_n1500_n27171# 0.0172f
C227 a_n1500_19797# w_n1594_21030# 0.0172f
C228 a_n1500_27213# a_n1500_25977# 3.11f
C229 a_n1500_28449# a_1500_28546# 0.217f
C230 a_n1500_n60543# a_1500_n60446# 0.217f
C231 w_n1594_n60546# a_1500_n59210# 0.0023f
C232 w_n1594_n63018# a_1500_n61682# 0.0023f
C233 a_n1500_n18519# a_n1500_n17283# 3.11f
C234 a_n1558_n6062# w_n1594_n7398# 0.0023f
C235 a_1500_29782# a_1500_28546# 0.0105f
C236 a_n1500_n11103# w_n1594_n9870# 0.0172f
C237 a_n1500_n2451# w_n1594_n2454# 1.65f
C238 a_n1558_12478# w_n1594_11142# 0.0023f
C239 a_n1500_16089# w_n1594_14850# 0.0172f
C240 a_1500_22366# a_1500_23602# 0.0105f
C241 w_n1594_n12342# a_n1500_n13575# 0.0172f
C242 w_n1594_n13578# a_n1558_n14714# 0.0023f
C243 w_n1594_3726# a_n1558_5062# 0.0023f
C244 a_n1500_38337# w_n1594_38334# 1.65f
C245 a_n1500_n54363# a_n1500_n55599# 3.11f
C246 a_n1500_45753# a_n1500_46989# 3.11f
C247 a_1500_52030# a_n1500_51933# 0.217f
C248 a_n1558_13714# w_n1594_12378# 0.0023f
C249 w_n1594_n34590# a_n1558_n33254# 0.0023f
C250 w_n1594_1254# a_n1500_2493# 0.0172f
C251 a_n1500_n20991# a_n1500_n22227# 3.11f
C252 a_n1558_n6062# w_n1594_n4926# 0.0023f
C253 a_1500_n40670# a_1500_n41906# 0.0105f
C254 a_n1500_n42003# a_n1558_n41906# 0.217f
C255 a_n1500_n49419# a_n1500_n50655# 3.11f
C256 a_n1500_n3687# w_n1594_n4926# 0.0172f
C257 a_n1500_30921# w_n1594_32154# 0.0172f
C258 w_n1594_32154# a_1500_31018# 0.0023f
C259 a_n1558_n15950# a_n1558_n14714# 0.0105f
C260 a_n1500_n16047# w_n1594_n14814# 0.0172f
C261 a_n1500_n34587# a_1500_n34490# 0.217f
C262 a_n1500_n18519# w_n1594_n18522# 1.65f
C263 a_n1500_n53127# w_n1594_n51894# 0.0172f
C264 w_n1594_38334# a_1500_37198# 0.0023f
C265 a_n1558_5062# a_n1558_3826# 0.0105f
C266 w_n1594_11142# a_n1500_11145# 1.65f
C267 w_n1594_38334# a_n1558_37198# 0.0023f
C268 a_n1500_n58071# a_1500_n57974# 0.217f
C269 w_n1594_18558# a_1500_18658# 0.0187f
C270 a_n1500_35865# a_n1500_34629# 3.11f
C271 w_n1594_18# a_n1558_n1118# 0.0023f
C272 a_n1558_35962# w_n1594_34626# 0.0023f
C273 a_n1500_n4923# a_1500_n4826# 0.217f
C274 a_1500_50794# w_n1594_49458# 0.0023f
C275 a_n1500_n23463# a_n1500_n24699# 3.11f
C276 a_n1500_n37059# w_n1594_n37062# 1.65f
C277 w_n1594_18# a_n1558_1354# 0.0023f
C278 a_1500_n32018# w_n1594_n32118# 0.0187f
C279 w_n1594_n56838# a_n1500_n56835# 1.65f
C280 a_n1558_39670# w_n1594_39570# 0.0187f
C281 a_n1558_n32018# w_n1594_n33354# 0.0023f
C282 a_n1500_45753# a_n1558_45850# 0.217f
C283 a_n1500_27213# w_n1594_27210# 1.65f
C284 a_n1500_n35823# a_1500_n35726# 0.217f
C285 w_n1594_n60546# a_n1500_n59307# 0.0172f
C286 w_n1594_n54366# a_n1500_n53127# 0.0172f
C287 w_n1594_55638# a_n1558_55738# 0.0187f
C288 a_n1500_29685# w_n1594_30918# 0.0172f
C289 w_n1594_n42006# a_n1500_n42003# 1.65f
C290 a_n1500_n29643# w_n1594_n29646# 1.65f
C291 a_1500_n9770# a_1500_n11006# 0.0105f
C292 w_n1594_1254# a_1500_1354# 0.0187f
C293 a_n1500_51933# a_n1500_50697# 3.11f
C294 a_n1500_3729# a_1500_3826# 0.217f
C295 a_1500_13714# w_n1594_13614# 0.0187f
C296 w_n1594_61818# a_n1500_60585# 0.0172f
C297 w_n1594_n58074# a_n1500_n58071# 1.65f
C298 a_n1500_46989# a_1500_47086# 0.217f
C299 a_n1500_17325# w_n1594_18558# 0.0172f
C300 a_n1500_n39531# a_n1558_n39434# 0.217f
C301 a_n1558_7534# w_n1594_7434# 0.0187f
C302 w_n1594_19794# a_1500_18658# 0.0023f
C303 a_1500_n11006# w_n1594_n9870# 0.0023f
C304 a_n1558_n11006# a_n1500_n11103# 0.217f
C305 a_n1500_n30879# a_1500_n30782# 0.217f
C306 a_n1558_31018# w_n1594_29682# 0.0023f
C307 a_n1558_12478# a_n1558_13714# 0.0105f
C308 a_1500_n45614# w_n1594_n46950# 0.0023f
C309 a_n1558_n8534# a_n1558_n9770# 0.0105f
C310 a_n1558_n59210# a_n1558_n60446# 0.0105f
C311 a_n1558_22366# w_n1594_21030# 0.0023f
C312 a_n1500_n39531# w_n1594_n38298# 0.0172f
C313 w_n1594_n2454# a_1500_n1118# 0.0023f
C314 w_n1594_n7398# a_1500_n8534# 0.0023f
C315 a_1500_44614# w_n1594_44514# 0.0187f
C316 a_n1500_n45711# a_n1558_n45614# 0.217f
C317 a_1500_n44378# a_1500_n45614# 0.0105f
C318 a_n1500_16089# a_1500_16186# 0.217f
C319 w_n1594_n43242# a_1500_n44378# 0.0023f
C320 a_n1558_17422# w_n1594_16086# 0.0023f
C321 w_n1594_8670# a_1500_10006# 0.0023f
C322 a_n1558_8770# a_n1500_8673# 0.217f
C323 a_n1500_30921# a_n1500_29685# 3.11f
C324 a_n1558_61918# a_n1558_60682# 0.0105f
C325 w_n1594_n59310# a_n1500_n60543# 0.0172f
C326 a_1500_42142# w_n1594_43278# 0.0023f
C327 a_1500_11242# w_n1594_11142# 0.0187f
C328 a_n1558_11242# w_n1594_12378# 0.0023f
C329 a_n1558_n36962# w_n1594_n35826# 0.0023f
C330 a_n1500_27213# w_n1594_28446# 0.0172f
C331 w_n1594_46986# a_n1500_46989# 1.65f
C332 a_1500_n24602# a_n1500_n24699# 0.217f
C333 a_1500_n23366# w_n1594_n22230# 0.0023f
C334 a_n1558_n33254# a_n1558_n34490# 0.0105f
C335 a_n1558_n15950# w_n1594_n14814# 0.0023f
C336 a_n1500_n2451# w_n1594_n3690# 0.0172f
C337 a_n1500_n18519# w_n1594_n17286# 0.0172f
C338 a_n1500_n51891# w_n1594_n51894# 1.65f
C339 a_n1558_22366# a_n1558_23602# 0.0105f
C340 a_n1558_8770# w_n1594_7434# 0.0023f
C341 w_n1594_n13578# a_n1500_n13575# 1.65f
C342 a_1500_n50558# w_n1594_n50658# 0.0187f
C343 a_n1558_n56738# a_n1558_n57974# 0.0105f
C344 a_n1558_40906# w_n1594_40806# 0.0187f
C345 a_1500_52030# w_n1594_50694# 0.0023f
C346 w_n1594_n30882# a_1500_n30782# 0.0187f
C347 w_n1594_54402# a_1500_53266# 0.0023f
C348 w_n1594_n45714# a_n1500_n44475# 0.0172f
C349 a_n1500_35865# a_n1558_35962# 0.217f
C350 a_n1500_n35823# w_n1594_n37062# 0.0172f
C351 a_n1500_9909# w_n1594_11142# 0.0172f
C352 a_n1500_40809# a_n1500_39573# 3.11f
C353 w_n1594_n56838# a_n1500_n55599# 0.0172f
C354 a_n1500_n59307# a_n1500_n60543# 3.11f
C355 w_n1594_59346# a_n1558_58210# 0.0023f
C356 w_n1594_60582# a_n1500_61821# 0.0172f
C357 a_n1558_45850# w_n1594_46986# 0.0023f
C358 a_n1558_35962# w_n1594_37098# 0.0023f
C359 a_n1500_33393# w_n1594_32154# 0.0172f
C360 w_n1594_n42006# a_n1500_n40767# 0.0172f
C361 a_1500_n43142# w_n1594_n44478# 0.0023f
C362 a_1500_n14714# a_1500_n15950# 0.0105f
C363 a_n1500_n1215# w_n1594_n2454# 0.0172f
C364 w_n1594_38334# a_n1558_39670# 0.0023f
C365 w_n1594_n58074# a_n1500_n56835# 0.0172f
C366 a_n1500_27213# w_n1594_25974# 0.0172f
C367 a_n1500_39573# w_n1594_39570# 1.65f
C368 a_n1558_52030# a_n1500_51933# 0.217f
C369 a_n1558_n17186# w_n1594_n16050# 0.0023f
C370 a_n1558_n29546# a_n1558_n30782# 0.0105f
C371 a_1500_34726# w_n1594_34626# 0.0187f
C372 a_n1500_n23463# w_n1594_n22230# 0.0172f
C373 a_n1558_56974# a_n1500_56877# 0.217f
C374 a_n1558_11242# a_n1558_12478# 0.0105f
C375 a_n1500_19797# w_n1594_18558# 0.0172f
C376 w_n1594_n34590# a_1500_n35726# 0.0023f
C377 a_1500_n11006# a_n1500_n11103# 0.217f
C378 a_n1500_n38295# w_n1594_n38298# 1.65f
C379 w_n1594_42042# a_n1500_43281# 0.0172f
C380 w_n1594_50694# a_n1500_50697# 1.65f
C381 a_n1558_34726# w_n1594_34626# 0.0187f
C382 w_n1594_13614# a_n1558_14950# 0.0023f
C383 a_1500_n19658# a_1500_n18422# 0.0105f
C384 a_n1558_7534# w_n1594_6198# 0.0023f
C385 a_n1558_24838# a_n1558_23602# 0.0105f
C386 a_1500_n9770# a_1500_n8534# 0.0105f
C387 a_n1500_n49419# w_n1594_n48186# 0.0172f
C388 a_n1500_n11103# a_n1500_n12339# 3.11f
C389 a_n1500_n53127# a_n1500_n54363# 3.11f
C390 a_1500_n61682# a_1500_n62918# 0.0105f
C391 a_n1500_n63015# a_n1558_n62918# 0.217f
C392 a_n1500_n50655# a_n1500_n51891# 3.11f
C393 w_n1594_n19758# a_n1500_n19755# 1.65f
C394 a_1500_n39434# a_1500_n40670# 0.0105f
C395 a_n1500_n40767# a_n1558_n40670# 0.217f
C396 a_1500_22366# w_n1594_22266# 0.0187f
C397 a_1500_11242# a_1500_10006# 0.0105f
C398 w_n1594_4962# a_n1500_4965# 1.65f
C399 a_n1558_11242# a_n1500_11145# 0.217f
C400 a_n1558_n35726# w_n1594_n35826# 0.0187f
C401 a_n1500_n48183# a_n1500_n49419# 3.11f
C402 a_n1558_31018# a_n1558_29782# 0.0105f
C403 a_n1558_n24602# a_n1558_n23366# 0.0105f
C404 w_n1594_n9870# a_1500_n8534# 0.0023f
C405 a_n1500_n33351# a_1500_n33254# 0.217f
C406 a_n1558_16186# w_n1594_16086# 0.0187f
C407 a_1500_43378# w_n1594_42042# 0.0023f
C408 w_n1594_29682# a_n1558_28546# 0.0023f
C409 a_n1500_29685# w_n1594_28446# 0.0172f
C410 a_n1500_n50655# w_n1594_n49422# 0.0172f
C411 a_n1500_n56835# a_1500_n56738# 0.217f
C412 a_1500_n49322# w_n1594_n50658# 0.0023f
C413 a_n1500_28449# a_n1500_27213# 3.11f
C414 a_1500_27310# a_1500_26074# 0.0105f
C415 w_n1594_19794# a_n1500_19797# 1.65f
C416 a_1500_n7298# a_1500_n8534# 0.0105f
C417 a_n1500_42045# w_n1594_42042# 1.65f
C418 a_1500_42142# w_n1594_40806# 0.0023f
C419 w_n1594_n1218# a_n1558_n1118# 0.0187f
C420 a_n1558_59446# a_n1558_58210# 0.0105f
C421 w_n1594_n30882# a_1500_n29546# 0.0023f
C422 a_n1558_18658# a_n1500_18561# 0.217f
C423 a_1500_n38198# a_1500_n39434# 0.0105f
C424 a_n1558_54502# w_n1594_55638# 0.0023f
C425 a_n1500_9909# a_1500_10006# 0.217f
C426 w_n1594_n55602# a_n1558_n56738# 0.0023f
C427 a_n1558_n32018# a_n1558_n30782# 0.0105f
C428 a_n1500_30921# w_n1594_29682# 0.0172f
C429 w_n1594_29682# a_1500_31018# 0.0023f
C430 a_n1500_14853# w_n1594_14850# 1.65f
C431 a_n1500_49461# a_n1558_49558# 0.217f
C432 a_n1558_n24602# a_n1558_n25838# 0.0105f
C433 a_n1500_38337# w_n1594_37098# 0.0172f
C434 a_n1500_n24699# w_n1594_n25938# 0.0172f
C435 a_n1500_23505# a_n1558_23602# 0.217f
C436 a_1500_n29546# w_n1594_n28410# 0.0023f
C437 a_n1558_16186# a_n1558_17422# 0.0105f
C438 a_n1558_21130# a_n1500_21033# 0.217f
C439 a_n1500_21# w_n1594_1254# 0.0172f
C440 a_1500_n9770# w_n1594_n11106# 0.0023f
C441 w_n1594_54402# a_n1558_55738# 0.0023f
C442 w_n1594_24738# a_n1558_23602# 0.0023f
C443 a_1500_8770# a_1500_10006# 0.0105f
C444 a_1500_n22130# w_n1594_n20994# 0.0023f
C445 a_1500_n36962# a_1500_n38198# 0.0105f
C446 a_n1500_n38295# a_n1558_n38198# 0.217f
C447 w_n1594_37098# a_1500_37198# 0.0187f
C448 a_n1558_44614# w_n1594_44514# 0.0187f
C449 a_n1500_n29643# a_1500_n29546# 0.217f
C450 w_n1594_37098# a_n1558_37198# 0.0187f
C451 a_n1500_n20991# a_n1500_n19755# 3.11f
C452 w_n1594_59346# a_1500_58210# 0.0023f
C453 a_n1500_12381# w_n1594_13614# 0.0172f
C454 w_n1594_44514# a_n1500_44517# 1.65f
C455 a_n1500_n46947# w_n1594_n45714# 0.0172f
C456 a_n1558_54502# a_n1558_55738# 0.0105f
C457 w_n1594_n16050# a_n1558_n14714# 0.0023f
C458 a_n1500_21033# w_n1594_22266# 0.0172f
C459 a_n1500_n37059# w_n1594_n38298# 0.0172f
C460 a_n1500_39573# w_n1594_38334# 0.0172f
C461 a_1500_38434# a_1500_39670# 0.0105f
C462 a_n1558_n4826# w_n1594_n4926# 0.0187f
C463 a_1500_n45614# w_n1594_n44478# 0.0023f
C464 a_n1500_n1215# a_n1558_n1118# 0.217f
C465 a_n1500_n25935# w_n1594_n27174# 0.0172f
C466 a_n1558_52030# w_n1594_50694# 0.0023f
C467 a_n1500_n48183# w_n1594_n48186# 1.65f
C468 a_1500_39670# w_n1594_39570# 0.0187f
C469 a_1500_34726# a_1500_33490# 0.0105f
C470 w_n1594_n30882# a_1500_n32018# 0.0023f
C471 w_n1594_44514# a_n1500_43281# 0.0172f
C472 a_1500_60682# a_1500_61918# 0.0105f
C473 a_1500_n6062# w_n1594_n6162# 0.0187f
C474 a_n1500_14853# a_n1500_13617# 3.11f
C475 w_n1594_49458# a_n1500_50697# 0.0172f
C476 a_1500_n8534# a_n1500_n8631# 0.217f
C477 a_1500_5062# a_n1500_4965# 0.217f
C478 w_n1594_4962# a_1500_3826# 0.0023f
C479 a_n1558_n8534# w_n1594_n7398# 0.0023f
C480 a_n1558_7534# w_n1594_8670# 0.0023f
C481 a_n1558_n32018# a_n1558_n33254# 0.0105f
C482 a_n1558_12478# w_n1594_13614# 0.0023f
C483 a_1500_33490# w_n1594_33390# 0.0187f
C484 a_n1558_2590# a_n1500_2493# 0.217f
C485 a_n1558_47086# a_n1558_48322# 0.0105f
C486 w_n1594_55638# a_1500_56974# 0.0023f
C487 a_n1500_n49419# w_n1594_n49422# 1.65f
C488 a_n1558_n55502# a_n1558_n56738# 0.0105f
C489 a_n1500_n6159# a_n1500_n7395# 3.11f
C490 a_n1500_49461# a_n1500_48225# 3.11f
C491 a_1500_32254# w_n1594_32154# 0.0187f
C492 a_1500_44614# a_n1500_44517# 0.217f
C493 w_n1594_n19758# a_1500_n20894# 0.0023f
C494 a_n1558_29782# w_n1594_30918# 0.0023f
C495 a_n1500_n43239# a_n1500_n44475# 3.11f
C496 a_1500_16186# w_n1594_17322# 0.0023f
C497 a_n1558_42142# w_n1594_43278# 0.0023f
C498 a_n1500_28449# a_n1500_29685# 3.11f
C499 a_1500_43378# w_n1594_44514# 0.0023f
C500 a_1500_n22130# w_n1594_n23466# 0.0023f
C501 w_n1594_18# a_n1558_118# 0.0187f
C502 w_n1594_n7398# a_n1558_n7298# 0.0187f
C503 a_n1500_33393# w_n1594_34626# 0.0172f
C504 a_n1500_40809# w_n1594_40806# 1.65f
C505 a_n1500_29685# a_1500_29782# 0.217f
C506 w_n1594_n8634# a_n1558_n9770# 0.0023f
C507 w_n1594_n55602# a_n1558_n55502# 0.0187f
C508 a_1500_n7298# w_n1594_n6162# 0.0023f
C509 a_n1558_14950# w_n1594_16086# 0.0023f
C510 a_n1500_3729# w_n1594_3726# 1.65f
C511 a_n1558_19894# a_n1558_18658# 0.0105f
C512 a_1500_n50558# w_n1594_n51894# 0.0023f
C513 w_n1594_n19758# a_n1558_n20894# 0.0023f
C514 w_n1594_58110# a_n1500_58113# 1.65f
C515 a_n1558_n11006# w_n1594_n11106# 0.0187f
C516 a_n1558_33490# w_n1594_33390# 0.0187f
C517 a_1500_n28310# w_n1594_n28410# 0.0187f
C518 a_n1558_33490# a_n1558_34726# 0.0105f
C519 a_n1500_14853# a_1500_14950# 0.217f
C520 a_n1558_29782# a_n1558_28546# 0.0105f
C521 a_n1558_8770# w_n1594_8670# 0.0187f
C522 a_n1558_n54266# w_n1594_n53130# 0.0023f
C523 a_1500_n23366# a_1500_n22130# 0.0105f
C524 w_n1594_n54366# a_1500_n55502# 0.0023f
C525 a_n1558_n28310# a_n1558_n29546# 0.0105f
C526 a_n1500_3729# a_n1558_3826# 0.217f
C527 a_n1500_n45711# w_n1594_n45714# 1.65f
C528 w_n1594_59346# a_n1500_59349# 1.65f
C529 a_1500_55738# w_n1594_56874# 0.0023f
C530 a_n1558_n41906# w_n1594_n40770# 0.0023f
C531 a_n1500_n19755# a_n1558_n19658# 0.217f
C532 a_n1500_59349# a_n1500_60585# 3.11f
C533 a_n1500_n11103# w_n1594_n11106# 1.65f
C534 w_n1594_n61782# a_n1558_n62918# 0.0023f
C535 w_n1594_n59310# a_n1558_n57974# 0.0023f
C536 a_n1500_n34587# a_n1500_n35823# 3.11f
C537 a_1500_43378# a_1500_44614# 0.0105f
C538 a_n1500_8673# w_n1594_7434# 0.0172f
C539 a_n1500_n25935# w_n1594_n25938# 1.65f
C540 a_1500_n44378# w_n1594_n44478# 0.0187f
C541 a_1500_24838# w_n1594_24738# 0.0187f
C542 a_n1500_n20991# a_1500_n20894# 0.217f
C543 a_n1558_n23366# w_n1594_n24702# 0.0023f
C544 a_n1500_n46947# w_n1594_n48186# 0.0172f
C545 w_n1594_n27174# a_1500_n27074# 0.0187f
C546 w_n1594_n28410# a_n1558_n27074# 0.0023f
C547 a_n1500_n51891# a_n1500_n53127# 3.11f
C548 w_n1594_8670# a_n1558_10006# 0.0023f
C549 a_n1500_38337# a_n1500_37101# 3.11f
C550 a_n1500_n17283# w_n1594_n18522# 0.0172f
C551 a_1500_n60446# a_1500_n61682# 0.0105f
C552 a_n1500_n61779# a_n1558_n61682# 0.217f
C553 a_n1558_1354# a_n1500_1257# 0.217f
C554 a_n1500_n16047# a_n1500_n14811# 3.11f
C555 a_1500_27310# a_1500_28546# 0.0105f
C556 w_n1594_n60546# a_n1558_n61682# 0.0023f
C557 a_n1558_n39434# w_n1594_n39534# 0.0187f
C558 a_n1500_49461# a_1500_49558# 0.217f
C559 w_n1594_n58074# a_n1558_n59210# 0.0023f
C560 a_n1558_n39434# w_n1594_n40770# 0.0023f
C561 a_n1500_n46947# a_n1500_n48183# 3.11f
C562 a_1500_3826# a_1500_5062# 0.0105f
C563 a_n1500_n20991# a_n1558_n20894# 0.217f
C564 a_1500_35962# a_1500_37198# 0.0105f
C565 a_n1500_n32115# a_1500_n32018# 0.217f
C566 a_n1558_n28310# a_n1500_n28407# 0.217f
C567 w_n1594_38334# a_1500_39670# 0.0023f
C568 a_1500_n28310# a_1500_n27074# 0.0105f
C569 w_n1594_55638# a_n1500_56877# 0.0172f
C570 a_n1500_37101# a_1500_37198# 0.217f
C571 a_1500_22366# a_n1500_22269# 0.217f
C572 w_n1594_59346# a_1500_59446# 0.0187f
C573 w_n1594_59346# a_1500_60682# 0.0023f
C574 w_n1594_n50658# a_1500_n51794# 0.0023f
C575 a_n1500_n18519# a_1500_n18422# 0.217f
C576 a_n1500_n48183# w_n1594_n49422# 0.0172f
C577 w_n1594_n2454# a_n1558_n2354# 0.0187f
C578 a_n1500_37101# a_n1558_37198# 0.217f
C579 a_n1500_n55599# a_1500_n55502# 0.217f
C580 a_n1558_5062# w_n1594_6198# 0.0023f
C581 a_1500_60682# a_n1500_60585# 0.217f
C582 a_1500_34726# a_1500_35962# 0.0105f
C583 a_n1558_n25838# w_n1594_n24702# 0.0023f
C584 a_n1500_n50655# a_1500_n50558# 0.217f
C585 w_n1594_45750# a_n1500_46989# 0.0172f
C586 a_n1500_18561# w_n1594_17322# 0.0172f
C587 a_n1558_n8534# w_n1594_n9870# 0.0023f
C588 a_1500_n14714# a_1500_n13478# 0.0105f
C589 w_n1594_n22230# a_n1500_n22227# 1.65f
C590 w_n1594_n55602# a_n1558_n54266# 0.0023f
C591 a_n1558_53266# w_n1594_53166# 0.0187f
C592 a_1500_17422# w_n1594_17322# 0.0187f
C593 w_n1594_60582# a_n1558_60682# 0.0187f
C594 w_n1594_55638# a_n1500_55641# 1.65f
C595 a_n1558_7534# a_n1558_6298# 0.0105f
C596 a_n1558_48322# a_n1558_49558# 0.0105f
C597 a_n1558_54502# w_n1594_54402# 0.0187f
C598 a_1500_n34490# w_n1594_n35826# 0.0023f
C599 a_n1558_42142# w_n1594_40806# 0.0023f
C600 a_1500_21130# w_n1594_22266# 0.0023f
C601 a_1500_n38198# w_n1594_n37062# 0.0023f
C602 a_1500_n24602# a_1500_n25838# 0.0105f
C603 a_n1500_59349# a_n1558_59446# 0.217f
C604 a_1500_n11006# w_n1594_n11106# 0.0187f
C605 a_1500_n19658# a_n1500_n19755# 0.217f
C606 a_n1500_n34587# w_n1594_n33354# 0.0172f
C607 w_n1594_n19758# a_n1500_n20991# 0.0172f
C608 a_n1558_n53030# w_n1594_n53130# 0.0187f
C609 a_n1500_n27171# a_n1500_n28407# 3.11f
C610 w_n1594_n17286# a_1500_n15950# 0.0023f
C611 w_n1594_n56838# a_1500_n57974# 0.0023f
C612 a_n1500_n37059# a_n1558_n36962# 0.217f
C613 a_1500_n35726# a_1500_n36962# 0.0105f
C614 w_n1594_n54366# a_1500_n54266# 0.0187f
C615 a_n1500_49461# w_n1594_50694# 0.0172f
C616 a_n1500_n45711# a_n1500_n44475# 3.11f
C617 a_n1500_33393# a_1500_33490# 0.217f
C618 a_n1500_28449# w_n1594_29682# 0.0172f
C619 w_n1594_50694# a_n1558_49558# 0.0023f
C620 a_n1500_18561# a_1500_18658# 0.217f
C621 a_n1558_45850# w_n1594_45750# 0.0187f
C622 w_n1594_n42006# a_1500_n43142# 0.0023f
C623 w_n1594_n43242# a_n1558_n43142# 0.0187f
C624 a_1500_n30782# w_n1594_n29646# 0.0023f
C625 a_n1500_n6159# a_n1500_n4923# 3.11f
C626 a_1500_29782# w_n1594_29682# 0.0187f
C627 w_n1594_53166# a_n1500_54405# 0.0172f
C628 a_n1558_n40670# w_n1594_n39534# 0.0023f
C629 w_n1594_n11106# a_n1500_n12339# 0.0172f
C630 a_n1558_n40670# w_n1594_n40770# 0.0187f
C631 a_n1500_55641# a_n1558_55738# 0.217f
C632 a_1500_18658# a_1500_17422# 0.0105f
C633 w_n1594_n61782# a_n1558_n61682# 0.0187f
C634 a_1500_39670# a_1500_40906# 0.0105f
C635 a_1500_55738# a_1500_54502# 0.0105f
C636 w_n1594_48222# a_1500_48322# 0.0187f
C637 w_n1594_23502# a_n1558_23602# 0.0187f
C638 a_n1500_21033# a_n1500_22269# 3.11f
C639 w_n1594_n13578# a_n1500_n14811# 0.0172f
C640 a_n1558_n30782# w_n1594_n32118# 0.0023f
C641 a_n1500_45753# w_n1594_44514# 0.0172f
C642 w_n1594_58110# a_1500_56974# 0.0023f
C643 a_n1558_n48086# w_n1594_n46950# 0.0023f
C644 a_n1558_29782# w_n1594_28446# 0.0023f
C645 w_n1594_n25938# a_1500_n27074# 0.0023f
C646 w_n1594_n27174# a_1500_n25838# 0.0023f
C647 a_n1500_n9867# a_n1558_n9770# 0.217f
C648 a_n1500_n17283# w_n1594_n17286# 1.65f
C649 a_n1558_16186# a_n1558_14950# 0.0105f
C650 w_n1594_n60546# a_n1558_n60446# 0.0187f
C651 a_n1558_24838# w_n1594_24738# 0.0187f
C652 a_n1558_n38198# w_n1594_n39534# 0.0023f
C653 w_n1594_n63018# a_n1558_n62918# 0.0187f
C654 a_n1500_33393# a_n1558_33490# 0.217f
C655 a_n1558_n22130# w_n1594_n22230# 0.0187f
C656 a_n1558_44614# a_n1500_44517# 0.217f
C657 a_n1500_16089# w_n1594_16086# 1.65f
C658 a_n1500_18561# a_n1500_17325# 3.11f
C659 a_n1558_n20894# a_n1558_n19658# 0.0105f
C660 a_n1558_n54266# a_n1558_n55502# 0.0105f
C661 a_n1500_48225# a_n1558_48322# 0.217f
C662 a_n1500_17325# a_1500_17422# 0.217f
C663 w_n1594_n34590# a_n1500_n34587# 1.65f
C664 a_n1500_n42003# a_n1500_n43239# 3.11f
C665 a_n1558_n49322# a_n1558_n50558# 0.0105f
C666 a_n1558_n24602# w_n1594_n24702# 0.0187f
C667 w_n1594_n1218# a_n1558_118# 0.0023f
C668 a_n1558_n8534# a_n1500_n8631# 0.217f
C669 a_n1558_27310# a_n1500_27213# 0.217f
C670 a_1500_n53030# w_n1594_n51894# 0.0023f
C671 w_n1594_n4926# a_1500_n4826# 0.0187f
C672 a_n1500_9909# a_n1558_10006# 0.217f
C673 a_n1558_24838# a_n1558_26074# 0.0105f
C674 a_n1500_44517# a_n1500_43281# 3.11f
C675 w_n1594_n3690# a_n1558_n2354# 0.0023f
C676 a_n1558_n17186# a_n1558_n18422# 0.0105f
C677 w_n1594_n14814# a_n1558_n14714# 0.0187f
C678 a_n1558_n11006# w_n1594_n12342# 0.0023f
C679 a_n1558_40906# a_n1500_40809# 0.217f
C680 a_1500_34726# a_n1500_34629# 0.217f
C681 a_1500_40906# w_n1594_40806# 0.0187f
C682 a_1500_n36962# w_n1594_n37062# 0.0187f
C683 a_n1558_n2354# a_n1558_n1118# 0.0105f
C684 a_1500_13714# w_n1594_12378# 0.0023f
C685 a_1500_n23366# w_n1594_n23466# 0.0187f
C686 w_n1594_24738# a_n1500_23505# 0.0172f
C687 a_n1500_34629# w_n1594_33390# 0.0172f
C688 a_n1558_n6062# w_n1594_n6162# 0.0187f
C689 w_n1594_n56838# a_1500_n56738# 0.0187f
C690 a_n1500_51933# w_n1594_50694# 0.0172f
C691 a_n1558_n33254# w_n1594_n32118# 0.0023f
C692 a_n1558_n51794# w_n1594_n53130# 0.0023f
C693 a_n1558_n12242# a_n1558_n11006# 0.0105f
C694 a_n1500_n33351# w_n1594_n33354# 1.65f
C695 a_n1558_53266# w_n1594_51930# 0.0023f
C696 a_n1558_34726# a_n1500_34629# 0.217f
C697 w_n1594_n54366# a_1500_n53030# 0.0023f
C698 w_n1594_n19758# a_n1558_n19658# 0.0187f
C699 w_n1594_n43242# a_n1558_n41906# 0.0023f
C700 a_1500_n29546# w_n1594_n29646# 0.0187f
C701 w_n1594_n42006# a_1500_n41906# 0.0187f
C702 a_n1558_40906# w_n1594_39570# 0.0023f
C703 w_n1594_n4926# a_n1558_n3590# 0.0023f
C704 w_n1594_3726# a_n1500_2493# 0.0172f
C705 w_n1594_2490# a_1500_3826# 0.0023f
C706 a_n1500_58113# a_n1500_56877# 3.11f
C707 w_n1594_n61782# a_n1558_n60446# 0.0023f
C708 a_1500_n19658# a_1500_n20894# 0.0105f
C709 a_n1500_n11103# w_n1594_n12342# 0.0172f
C710 a_n1500_49461# w_n1594_49458# 1.65f
C711 w_n1594_n58074# a_1500_n57974# 0.0187f
C712 a_n1558_47086# w_n1594_46986# 0.0187f
C713 a_n1558_18658# a_n1558_17422# 0.0105f
C714 w_n1594_49458# a_n1558_49558# 0.0187f
C715 w_n1594_56874# a_n1558_58210# 0.0023f
C716 w_n1594_58110# a_n1500_56877# 0.0172f
C717 a_n1558_2590# w_n1594_2490# 0.0187f
C718 a_n1558_n46850# w_n1594_n46950# 0.0187f
C719 w_n1594_n25938# a_1500_n25838# 0.0187f
C720 a_1500_n59210# a_1500_n60446# 0.0105f
C721 a_n1500_n60543# a_n1558_n60446# 0.217f
C722 a_n1558_43378# a_n1558_42142# 0.0105f
C723 w_n1594_n63018# a_n1558_n61682# 0.0023f
C724 w_n1594_n60546# a_n1558_n59210# 0.0023f
C725 a_1500_n11006# a_1500_n12242# 0.0105f
C726 a_1500_43378# a_n1500_43281# 0.217f
C727 a_n1500_n45711# a_n1500_n46947# 3.11f
C728 a_n1558_26074# w_n1594_24738# 0.0023f
C729 a_n1500_14853# w_n1594_13614# 0.0172f
C730 a_n1558_31018# w_n1594_30918# 0.0187f
C731 w_n1594_4962# a_n1558_3826# 0.0023f
C732 a_1500_24838# w_n1594_23502# 0.0023f
C733 a_n1500_n23463# w_n1594_n23466# 1.65f
C734 a_n1500_32157# w_n1594_30918# 0.0172f
C735 a_n1500_n12339# a_1500_n12242# 0.217f
C736 a_n1500_n54363# a_1500_n54266# 0.217f
C737 a_n1500_42045# a_n1500_43281# 3.11f
C738 a_1500_2590# a_n1500_2493# 0.217f
C739 w_n1594_n34590# a_n1500_n33351# 0.0172f
C740 a_n1558_50794# w_n1594_51930# 0.0023f
C741 a_n1558_n4826# a_n1558_n6062# 0.0105f
C742 a_1500_n6062# a_1500_n4826# 0.0105f
C743 a_1500_49558# w_n1594_50694# 0.0023f
C744 w_n1594_n59310# a_1500_n60446# 0.0023f
C745 a_n1500_18561# a_n1500_19797# 3.11f
C746 a_n1500_n49419# a_1500_n49322# 0.217f
C747 w_n1594_n19758# a_n1558_n18422# 0.0023f
C748 w_n1594_61818# a_1500_60682# 0.0023f
C749 a_1500_n33254# a_1500_n34490# 0.0105f
C750 a_1500_n2354# w_n1594_n2454# 0.0187f
C751 a_n1500_n34587# a_n1558_n34490# 0.217f
C752 w_n1594_8670# a_n1500_8673# 1.65f
C753 a_1500_n51794# w_n1594_n51894# 0.0187f
C754 w_n1594_53166# a_1500_54502# 0.0023f
C755 a_n1558_35962# a_n1558_37198# 0.0105f
C756 a_n1500_6201# w_n1594_7434# 0.0172f
C757 a_n1558_19894# w_n1594_21030# 0.0023f
C758 a_n1500_n58071# a_n1558_n57974# 0.217f
C759 a_1500_n56738# a_1500_n57974# 0.0105f
C760 a_1500_32254# a_1500_33490# 0.0105f
C761 a_1500_27310# a_n1500_27213# 0.217f
C762 w_n1594_n19758# a_1500_n19658# 0.0187f
C763 w_n1594_54402# a_n1500_55641# 0.0172f
C764 a_1500_n35726# w_n1594_n37062# 0.0023f
C765 a_1500_24838# a_1500_23602# 0.0105f
C766 a_n1558_n3590# a_n1558_n2354# 0.0105f
C767 a_n1500_n23463# a_1500_n23366# 0.217f
C768 a_1500_45850# w_n1594_44514# 0.0023f
C769 a_n1558_22366# w_n1594_23502# 0.0023f
C770 a_1500_n11006# w_n1594_n12342# 0.0023f
C771 a_1500_n14714# w_n1594_n13578# 0.0023f
C772 a_n1500_32157# w_n1594_33390# 0.0172f
C773 a_n1558_n32018# w_n1594_n32118# 0.0187f
C774 w_n1594_n56838# a_1500_n55502# 0.0023f
C775 a_n1500_n32115# w_n1594_n33354# 0.0172f
C776 a_n1558_40906# a_n1558_42142# 0.0105f
C777 a_n1500_n35823# a_n1558_n35726# 0.217f
C778 w_n1594_48222# a_n1500_46989# 0.0172f
C779 w_n1594_49458# a_n1500_48225# 0.0172f
C780 a_n1500_30921# a_n1558_31018# 0.217f
C781 a_n1558_16186# a_n1500_16089# 0.217f
C782 w_n1594_n14814# a_n1500_n13575# 0.0172f
C783 a_n1558_38434# w_n1594_39570# 0.0023f
C784 a_1500_n28310# w_n1594_n29646# 0.0023f
C785 a_n1558_35962# a_n1558_34726# 0.0105f
C786 w_n1594_n42006# a_1500_n40670# 0.0023f
C787 a_n1500_30921# a_n1500_32157# 3.11f
C788 w_n1594_n12342# a_n1500_n12339# 1.65f
C789 a_1500_2590# a_1500_1354# 0.0105f
C790 a_n1558_21130# w_n1594_21030# 0.0187f
C791 a_n1558_5062# a_n1558_6298# 0.0105f
C792 a_1500_n9770# w_n1594_n8634# 0.0023f
C793 w_n1594_n58074# a_1500_n56738# 0.0023f
C794 a_n1500_n3687# w_n1594_n2454# 0.0172f
C795 a_1500_12478# w_n1594_11142# 0.0023f
C796 a_n1500_n18519# a_n1500_n19755# 3.11f
C797 w_n1594_3726# a_1500_5062# 0.0023f
C798 a_n1500_n30879# a_n1558_n30782# 0.217f
C799 a_1500_n29546# a_1500_n30782# 0.0105f
C800 a_n1558_n12242# a_n1500_n12339# 0.217f
C801 a_n1558_n6062# a_n1558_n7298# 0.0105f
C802 a_n1500_25977# w_n1594_24738# 0.0172f
C803 a_1500_n22130# a_n1500_n22227# 0.217f
C804 a_n1558_n45614# w_n1594_n46950# 0.0023f
C805 a_1500_n24602# w_n1594_n23466# 0.0023f
C806 a_1500_24838# w_n1594_25974# 0.0023f
C807 a_1500_n38198# w_n1594_n38298# 0.0187f
C808 a_1500_n3590# w_n1594_n4926# 0.0023f
C809 a_n1500_35865# w_n1594_35862# 1.65f
C810 a_1500_n7298# w_n1594_n8634# 0.0023f
C811 w_n1594_n43242# a_n1558_n44378# 0.0023f
C812 a_1500_45850# a_1500_44614# 0.0105f
C813 a_n1500_33393# a_n1500_34629# 3.11f
C814 w_n1594_56874# a_1500_58210# 0.0023f
C815 a_n1558_7534# a_n1500_7437# 0.217f
C816 a_1500_n49322# w_n1594_n48186# 0.0023f
C817 a_n1500_n16047# a_1500_n15950# 0.217f
C818 a_n1558_2590# w_n1594_1254# 0.0023f
C819 a_n1558_n53030# a_n1558_n54266# 0.0105f
C820 a_n1558_32254# w_n1594_32154# 0.0187f
C821 a_n1558_n50558# a_n1558_n51794# 0.0105f
C822 w_n1594_18# a_1500_n1118# 0.0023f
C823 a_1500_56974# a_n1500_56877# 0.217f
C824 w_n1594_n59310# a_1500_n59210# 0.0187f
C825 a_n1500_n40767# a_n1500_n42003# 3.11f
C826 a_n1558_n48086# a_n1558_n49322# 0.0105f
C827 a_n1500_n37059# w_n1594_n35826# 0.0172f
C828 a_n1558_n24602# a_n1500_n24699# 0.217f
C829 a_1500_n24602# a_1500_n23366# 0.0105f
C830 a_n1558_n23366# w_n1594_n22230# 0.0023f
C831 a_n1558_24838# w_n1594_23502# 0.0023f
C832 a_n1500_18561# w_n1594_18558# 1.65f
C833 w_n1594_2490# a_n1558_1354# 0.0023f
C834 a_n1558_26074# a_n1500_25977# 0.217f
C835 a_1500_50794# w_n1594_51930# 0.0023f
C836 a_n1558_19894# a_n1500_19797# 0.217f
C837 w_n1594_22266# a_n1558_23602# 0.0023f
C838 a_n1500_45753# a_n1500_44517# 3.11f
C839 w_n1594_9906# a_1500_10006# 0.0187f
C840 w_n1594_18558# a_1500_17422# 0.0023f
C841 a_1500_n50558# w_n1594_n49422# 0.0023f
C842 a_n1558_n50558# w_n1594_n50658# 0.0187f
C843 a_1500_49558# w_n1594_49458# 0.0187f
C844 a_n1500_61821# a_1500_61918# 0.217f
C845 w_n1594_n30882# a_n1558_n30782# 0.0187f
C846 a_1500_n17186# a_1500_n15950# 0.0105f
C847 a_n1500_n7395# w_n1594_n7398# 1.65f
C848 a_n1500_n39531# a_n1500_n40767# 3.11f
C849 a_1500_n2354# w_n1594_n3690# 0.0023f
C850 w_n1594_61818# a_n1558_61918# 0.0187f
C851 a_n1500_n16047# a_n1500_n17283# 3.11f
C852 a_1500_n32018# a_1500_n30782# 0.0105f
C853 w_n1594_53166# a_n1500_53169# 1.65f
C854 a_n1500_6201# w_n1594_6198# 1.65f
C855 a_n1500_n59307# a_1500_n59210# 0.217f
C856 w_n1594_60582# a_1500_61918# 0.0023f
C857 a_n1500_12381# w_n1594_12378# 1.65f
C858 w_n1594_7434# a_1500_6298# 0.0023f
C859 a_n1500_14853# w_n1594_16086# 0.0172f
C860 w_n1594_n16050# a_n1500_n14811# 0.0172f
C861 a_n1500_n25935# a_n1558_n25838# 0.217f
C862 a_1500_n39434# w_n1594_n38298# 0.0023f
C863 a_n1558_n43142# w_n1594_n44478# 0.0023f
C864 a_n1500_9909# a_n1500_8673# 3.11f
C865 a_n1500_18561# w_n1594_19794# 0.0172f
C866 w_n1594_49458# a_n1558_48322# 0.0023f
C867 a_n1500_40809# w_n1594_39570# 0.0172f
C868 w_n1594_7434# a_n1558_6298# 0.0023f
C869 a_n1500_n38295# a_n1500_n39531# 3.11f
C870 a_1500_44614# w_n1594_43278# 0.0023f
C871 w_n1594_23502# a_n1500_23505# 1.65f
C872 a_n1558_17422# w_n1594_17322# 0.0187f
C873 a_n1558_38434# w_n1594_38334# 0.0187f
C874 w_n1594_n59310# a_n1500_n59307# 1.65f
C875 a_n1500_30921# w_n1594_30918# 1.65f
C876 w_n1594_n8634# a_n1500_n8631# 1.65f
C877 w_n1594_30918# a_1500_31018# 0.0187f
C878 a_1500_n17186# a_n1500_n17283# 0.217f
C879 a_n1558_26074# w_n1594_27210# 0.0023f
C880 a_1500_n46850# w_n1594_n45714# 0.0023f
C881 w_n1594_4962# a_n1558_5062# 0.0187f
C882 w_n1594_46986# a_n1500_48225# 0.0172f
C883 a_1500_8770# a_n1500_8673# 0.217f
C884 a_n1500_n1215# w_n1594_18# 0.0172f
C885 a_n1500_54405# a_1500_54502# 0.217f
C886 w_n1594_n13578# a_n1500_n12339# 0.0172f
C887 a_1500_38434# w_n1594_39570# 0.0023f
C888 a_1500_n36962# w_n1594_n38298# 0.0023f
C889 w_n1594_n34590# a_n1558_n35726# 0.0023f
C890 a_1500_34726# w_n1594_33390# 0.0023f
C891 w_n1594_n11106# a_1500_n12242# 0.0023f
C892 a_n1558_n18422# a_n1558_n19658# 0.0105f
C893 a_n1500_n3687# w_n1594_n3690# 1.65f
C894 a_n1558_12478# w_n1594_12378# 0.0187f
C895 a_n1558_24838# w_n1594_25974# 0.0023f
C896 a_n1500_33393# a_n1500_32157# 3.11f
C897 a_1500_8770# w_n1594_7434# 0.0023f
C898 a_1500_n48086# w_n1594_n48186# 0.0187f
C899 w_n1594_n20994# a_n1500_n22227# 0.0172f
C900 a_1500_n17186# w_n1594_n18522# 0.0023f
C901 a_n1500_n53127# a_1500_n53030# 0.217f
C902 a_n1558_34726# w_n1594_33390# 0.0023f
C903 a_1500_23602# a_n1500_23505# 0.217f
C904 a_1500_52030# w_n1594_53166# 0.0023f
C905 a_n1558_11242# w_n1594_9906# 0.0023f
C906 a_1500_n20894# w_n1594_n22230# 0.0023f
C907 a_n1500_n2451# w_n1594_n1218# 0.0172f
C908 a_n1500_n35823# w_n1594_n35826# 1.65f
C909 a_n1500_n48183# a_1500_n48086# 0.217f
C910 a_n1500_n33351# a_n1558_n33254# 0.217f
C911 a_1500_n32018# a_1500_n33254# 0.0105f
C912 a_n1500_17325# w_n1594_16086# 0.0172f
C913 w_n1594_n18522# a_1500_n18422# 0.0187f
C914 a_1500_23602# w_n1594_24738# 0.0023f
C915 a_n1500_13617# w_n1594_14850# 0.0172f
C916 a_n1558_12478# a_n1500_12381# 0.217f
C917 a_n1558_n4826# w_n1594_n6162# 0.0023f
C918 w_n1594_12378# a_n1500_11145# 0.0172f
C919 w_n1594_n22230# a_n1558_n20894# 0.0023f
C920 a_1500_n49322# w_n1594_n49422# 0.0187f
C921 a_n1558_19894# w_n1594_18558# 0.0023f
C922 a_n1500_30921# a_1500_31018# 0.217f
C923 a_1500_n55502# a_1500_n56738# 0.0105f
C924 a_n1558_n49322# w_n1594_n50658# 0.0023f
C925 a_n1500_n56835# a_n1558_n56738# 0.217f
C926 a_1500_n9770# a_n1500_n9867# 0.217f
C927 a_n1558_n13478# w_n1594_n12342# 0.0023f
C928 a_n1500_55641# a_n1500_56877# 3.11f
C929 a_1500_59446# a_1500_58210# 0.0105f
C930 w_n1594_n30882# a_n1558_n29546# 0.0023f
C931 a_n1500_n9867# w_n1594_n9870# 1.65f
C932 w_n1594_1254# a_n1558_1354# 0.0187f
C933 w_n1594_n55602# a_n1500_n56835# 0.0172f
C934 a_1500_42142# a_1500_40906# 0.0105f
C935 a_n1558_n13478# a_n1558_n12242# 0.0105f
C936 w_n1594_35862# a_1500_35962# 0.0187f
C937 a_n1500_12381# a_n1500_11145# 3.11f
C938 a_n1558_28546# w_n1594_27210# 0.0023f
C939 a_n1500_17325# a_n1558_17422# 0.217f
C940 a_n1558_n29546# w_n1594_n28410# 0.0023f
C941 a_n1558_56974# a_n1558_58210# 0.0105f
C942 a_n1558_n12242# w_n1594_n11106# 0.0023f
C943 a_n1500_61821# a_n1500_60585# 3.11f
C944 a_n1500_37101# w_n1594_35862# 0.0172f
C945 w_n1594_18# a_1500_118# 0.0187f
C946 a_n1500_25977# w_n1594_27210# 0.0172f
C947 w_n1594_14850# a_1500_16186# 0.0023f
C948 a_n1558_22366# a_n1558_21130# 0.0105f
C949 w_n1594_n19758# a_n1500_n18519# 0.0172f
C950 a_n1500_n16047# w_n1594_n17286# 0.0172f
C951 a_n1558_53266# a_n1500_53169# 0.217f
C952 w_n1594_51930# a_n1500_53169# 0.0172f
C953 a_n1558_n22130# w_n1594_n20994# 0.0023f
C954 w_n1594_2490# a_n1558_3826# 0.0023f
C955 a_n1558_19894# w_n1594_19794# 0.0187f
C956 a_n1558_43378# w_n1594_42042# 0.0023f
C957 w_n1594_n23466# a_n1500_n22227# 0.0172f
C958 w_n1594_14850# a_1500_14950# 0.0187f
C959 a_n1500_n1215# a_n1500_n2451# 3.11f
C960 a_1500_n28310# a_1500_n29546# 0.0105f
C961 w_n1594_6198# a_1500_6298# 0.0187f
C962 w_n1594_60582# a_n1500_60585# 1.65f
C963 a_n1500_n29643# a_n1558_n29546# 0.217f
C964 a_1500_n45614# w_n1594_n45714# 0.0187f
C965 a_1500_n7298# a_n1500_n7395# 0.217f
C966 a_1500_55738# w_n1594_55638# 0.0187f
C967 a_1500_22366# a_1500_21130# 0.0105f
C968 w_n1594_18# a_n1500_1257# 0.0172f
C969 a_n1558_22366# w_n1594_22266# 0.0187f
C970 w_n1594_46986# a_n1558_48322# 0.0023f
C971 a_1500_2590# w_n1594_2490# 0.0187f
C972 w_n1594_n6162# a_n1558_n7298# 0.0023f
C973 a_n1558_13714# w_n1594_14850# 0.0023f
C974 a_n1558_47086# w_n1594_45750# 0.0023f
C975 a_1500_n13478# a_1500_n12242# 0.0105f
C976 w_n1594_6198# a_n1558_6298# 0.0187f
C977 a_n1558_16186# w_n1594_17322# 0.0023f
C978 a_n1558_n34490# a_n1558_n35726# 0.0105f
C979 w_n1594_21030# a_n1500_22269# 0.0172f
C980 a_n1558_n45614# w_n1594_n44478# 0.0023f
C981 a_n1500_n24699# w_n1594_n24702# 1.65f
C982 w_n1594_29682# a_1500_28546# 0.0023f
C983 a_n1558_26074# w_n1594_25974# 0.0187f
C984 w_n1594_38334# a_1500_38434# 0.0187f
C985 w_n1594_n28410# a_n1500_n28407# 1.65f
C986 a_1500_n46850# w_n1594_n48186# 0.0023f
C987 a_n1500_n3687# a_n1558_n3590# 0.217f
C988 a_n1500_54405# a_n1500_53169# 3.11f
C989 a_1500_n17186# w_n1594_n17286# 0.0187f
C990 a_n1500_n4923# w_n1594_n4926# 1.65f
C991 a_n1558_n51794# a_n1558_n53030# 0.0105f
C992 a_n1558_21130# w_n1594_19794# 0.0023f
C993 w_n1594_n30882# a_n1558_n32018# 0.0023f
C994 w_n1594_n1218# a_1500_n1118# 0.0187f
C995 a_n1500_n61779# a_n1500_n63015# 3.11f
C996 a_1500_11242# w_n1594_12378# 0.0023f
C997 a_n1558_n46850# a_n1558_n48086# 0.0105f
C998 w_n1594_n17286# a_1500_n18422# 0.0023f
C999 a_n1500_n29643# a_n1500_n28407# 3.11f
C1000 w_n1594_28446# a_n1558_28546# 0.0187f
C1001 a_n1558_n14714# a_n1500_n14811# 0.217f
C1002 a_1500_n14714# w_n1594_n16050# 0.0023f
C1003 a_1500_n48086# w_n1594_n49422# 0.0023f
C1004 a_1500_7534# w_n1594_7434# 0.0187f
C1005 a_n1558_40906# w_n1594_42042# 0.0023f
C1006 a_n1500_n43239# a_1500_n43142# 0.217f
C1007 a_1500_52030# w_n1594_51930# 0.0187f
C1008 a_n1500_59349# a_1500_59446# 0.217f
C1009 a_n1558_n22130# w_n1594_n23466# 0.0023f
C1010 a_n1500_n9867# a_n1500_n8631# 3.11f
C1011 a_1500_53266# w_n1594_53166# 0.0187f
C1012 w_n1594_n55602# a_n1500_n55599# 1.65f
C1013 a_1500_n13478# w_n1594_n12342# 0.0023f
C1014 a_n1500_n20991# w_n1594_n22230# 0.0172f
C1015 a_n1558_n50558# w_n1594_n51894# 0.0023f
C1016 a_n1500_13617# a_n1558_13714# 0.217f
C1017 a_n1500_n6159# w_n1594_n7398# 0.0172f
C1018 w_n1594_11142# a_1500_10006# 0.0023f
C1019 w_n1594_59346# a_n1500_58113# 0.0172f
C1020 a_n1558_44614# w_n1594_43278# 0.0023f
C1021 w_n1594_60582# a_n1558_59446# 0.0023f
C1022 a_n1500_40809# a_1500_40906# 0.217f
C1023 a_n1500_33393# w_n1594_33390# 1.65f
C1024 a_n1500_n11103# a_n1500_n9867# 3.11f
C1025 w_n1594_43278# a_n1500_44517# 0.0172f
C1026 a_n1558_n28310# w_n1594_n28410# 0.0187f
C1027 a_1500_n28310# w_n1594_n27174# 0.0023f
C1028 a_n1558_n13478# w_n1594_n13578# 0.0187f
C1029 a_1500_21130# a_n1500_21033# 0.217f
C1030 a_n1500_n25935# a_n1500_n27171# 3.11f
C1031 a_n1500_n7395# a_n1500_n8631# 3.11f
C1032 a_1500_44614# w_n1594_45750# 0.0023f
C1033 a_n1500_n23463# a_n1500_n22227# 3.11f
C1034 a_n1500_n54363# w_n1594_n53130# 0.0172f
C1035 a_1500_n34490# w_n1594_n33354# 0.0023f
C1036 a_n1558_n59210# a_n1558_n57974# 0.0105f
C1037 a_n1500_n6159# w_n1594_n4926# 0.0172f
C1038 w_n1594_35862# a_n1500_34629# 0.0172f
C1039 a_n1558_n15950# w_n1594_n17286# 0.0023f
C1040 a_n1500_n37059# a_n1500_n38295# 3.11f
C1041 w_n1594_n54366# a_n1558_n55502# 0.0023f
C1042 a_n1500_n1215# a_1500_n1118# 0.217f
C1043 a_n1558_52030# w_n1594_53166# 0.0023f
C1044 a_1500_14950# a_1500_16186# 0.0105f
C1045 a_1500_32254# a_n1500_32157# 0.217f
C1046 a_1500_n44378# w_n1594_n45714# 0.0023f
C1047 a_n1500_21# a_n1558_118# 0.217f
C1048 w_n1594_n43242# a_n1500_n44475# 0.0172f
C1049 a_n1500_6201# a_1500_6298# 0.217f
C1050 a_1500_n2354# a_1500_n3590# 0.0105f
C1051 a_n1500_n1215# w_n1594_n1218# 1.65f
C1052 a_1500_40906# w_n1594_39570# 0.0023f
C1053 a_n1500_n42003# w_n1594_n40770# 0.0172f
C1054 a_n1500_38337# a_n1500_39573# 3.11f
C1055 a_1500_60682# a_1500_59446# 0.0105f
C1056 a_n1500_25977# w_n1594_25974# 1.65f
C1057 w_n1594_18# a_1500_1354# 0.0023f
C1058 a_n1558_8770# w_n1594_9906# 0.0023f
C1059 w_n1594_n61782# a_n1500_n63015# 0.0172f
C1060 w_n1594_43278# a_n1500_43281# 1.65f
C1061 a_n1558_43378# w_n1594_44514# 0.0023f
C1062 w_n1594_51930# a_n1500_50697# 0.0172f
C1063 w_n1594_n12342# a_1500_n12242# 0.0187f
C1064 w_n1594_n59310# a_n1500_n58071# 0.0172f
C1065 a_1500_12478# w_n1594_13614# 0.0023f
C1066 w_n1594_56874# a_n1558_56974# 0.0187f
C1067 a_n1558_n44378# w_n1594_n44478# 0.0187f
C1068 a_1500_n24602# w_n1594_n25938# 0.0023f
C1069 a_n1558_n8534# a_n1558_n7298# 0.0105f
C1070 a_n1500_6201# a_n1558_6298# 0.217f
C1071 w_n1594_n27174# a_n1558_n27074# 0.0187f
C1072 w_n1594_n28410# a_n1500_n27171# 0.0172f
C1073 a_n1500_n51891# a_1500_n51794# 0.217f
C1074 a_1500_26074# a_1500_24838# 0.0105f
C1075 a_1500_29782# w_n1594_30918# 0.0023f
C1076 a_n1500_n39531# w_n1594_n39534# 1.65f
C1077 w_n1594_n60546# a_n1500_n61779# 0.0172f
C1078 a_1500_11242# a_n1500_11145# 0.217f
C1079 a_n1500_n39531# w_n1594_n40770# 0.0172f
C1080 a_n1500_n46947# a_1500_n46850# 0.217f
C1081 w_n1594_n8634# a_1500_n8534# 0.0187f
C1082 a_1500_2590# w_n1594_1254# 0.0023f
C1083 a_n1500_n32115# a_n1558_n32018# 0.217f
C1084 a_1500_43378# w_n1594_43278# 0.0187f
C1085 a_n1500_9909# w_n1594_8670# 0.0172f
C1086 w_n1594_22266# a_n1500_23505# 0.0172f
C1087 a_n1558_38434# w_n1594_37098# 0.0023f
C1088 w_n1594_n50658# a_n1558_n51794# 0.0023f
C1089 a_n1500_7437# a_n1500_8673# 3.11f
C1090 w_n1594_n14814# a_n1500_n14811# 1.65f
C1091 a_n1500_n55599# a_n1558_n55502# 0.217f
C1092 w_n1594_9906# a_n1558_10006# 0.0187f
C1093 a_1500_n54266# a_1500_n55502# 0.0105f
C1094 a_n1500_n59307# a_n1500_n58071# 3.11f
C1095 w_n1594_n34590# a_1500_n34490# 0.0187f
C1096 a_n1500_42045# w_n1594_43278# 0.0172f
C1097 a_1500_n3590# a_n1500_n3687# 0.217f
C1098 a_n1558_n41906# a_n1558_n43142# 0.0105f
C1099 a_n1500_28449# a_n1558_28546# 0.217f
C1100 a_1500_42142# w_n1594_42042# 0.0187f
C1101 a_n1500_n50655# a_n1558_n50558# 0.217f
C1102 a_n1558_11242# w_n1594_11142# 0.0187f
C1103 a_1500_n49322# a_1500_n50558# 0.0105f
C1104 a_n1500_n25935# w_n1594_n24702# 0.0172f
C1105 a_n1500_14853# a_n1558_14950# 0.217f
C1106 a_n1500_7437# w_n1594_7434# 1.65f
C1107 a_n1500_9909# a_n1500_11145# 3.11f
C1108 a_1500_8770# w_n1594_8670# 0.0187f
C1109 w_n1594_n55602# a_n1500_n54363# 0.0172f
C1110 a_1500_23602# w_n1594_23502# 0.0187f
C1111 a_n1500_n13575# a_n1500_n14811# 3.11f
C1112 w_n1594_58110# a_n1558_59446# 0.0023f
C1113 a_n1500_n6159# a_1500_n6062# 0.217f
C1114 a_1500_n1118# a_1500_118# 0.0105f
C1115 a_1500_7534# w_n1594_6198# 0.0023f
C1116 a_n1500_45753# w_n1594_46986# 0.0172f
C1117 a_n1558_50794# a_n1500_50697# 0.217f
C1118 a_n1558_n34490# w_n1594_n35826# 0.0023f
C1119 a_n1558_n12242# w_n1594_n12342# 0.0187f
C1120 a_n1558_n38198# w_n1594_n37062# 0.0023f
C1121 w_n1594_n1218# a_1500_118# 0.0023f
C1122 a_n1558_33490# a_n1558_32254# 0.0105f
C1123 a_1500_n22130# a_1500_n20894# 0.0105f
C1124 a_1500_29782# a_1500_31018# 0.0105f
C1125 a_n1500_n53127# w_n1594_n53130# 1.65f
C1126 a_1500_53266# w_n1594_51930# 0.0023f
C1127 w_n1594_61818# a_n1500_61821# 1.65f
C1128 w_n1594_n56838# a_n1558_n57974# 0.0023f
C1129 a_n1500_n27171# a_1500_n27074# 0.217f
C1130 a_1500_n33254# w_n1594_n33354# 0.0187f
C1131 a_n1500_n19755# w_n1594_n20994# 0.0172f
C1132 w_n1594_n16050# a_1500_n15950# 0.0187f
C1133 a_1500_n13478# w_n1594_n13578# 0.0187f
C1134 a_n1558_n4826# w_n1594_n3690# 0.0023f
C1135 w_n1594_n54366# a_n1558_n54266# 0.0187f
C1136 a_1500_17422# a_1500_16186# 0.0105f
C1137 w_n1594_18558# a_n1558_17422# 0.0023f
C1138 a_1500_n44378# a_n1500_n44475# 0.217f
C1139 a_n1558_35962# w_n1594_35862# 0.0187f
C1140 w_n1594_n42006# a_n1558_n43142# 0.0023f
C1141 w_n1594_n43242# a_n1500_n43239# 1.65f
C1142 a_n1558_n30782# w_n1594_n29646# 0.0023f
C1143 a_n1500_n40767# w_n1594_n39534# 0.0172f
C1144 w_n1594_n6162# a_1500_n4826# 0.0023f
C1145 a_n1500_n40767# w_n1594_n40770# 1.65f
C1146 w_n1594_n61782# a_n1500_n61779# 1.65f
C1147 a_n1500_n19755# w_n1594_n18522# 0.0172f
C1148 a_1500_55738# w_n1594_54402# 0.0023f
C1149 a_1500_32254# w_n1594_30918# 0.0023f
C1150 a_n1500_n30879# w_n1594_n32118# 0.0172f
C1151 a_n1558_52030# w_n1594_51930# 0.0187f
C1152 a_n1558_52030# a_n1558_53266# 0.0105f
C1153 a_n1558_22366# a_n1500_22269# 0.217f
C1154 a_n1500_n48183# w_n1594_n46950# 0.0172f
C1155 a_n1500_n18519# a_n1558_n18422# 0.217f
C1156 w_n1594_n25938# a_n1558_n27074# 0.0023f
C1157 a_n1500_28449# w_n1594_27210# 0.0172f
C1158 a_1500_50794# a_1500_52030# 0.0105f
C1159 a_n1500_45753# a_1500_45850# 0.217f
C1160 a_1500_5062# w_n1594_6198# 0.0023f
C1161 a_n1500_n17283# w_n1594_n16050# 0.0172f
C1162 a_n1500_n38295# w_n1594_n39534# 0.0172f
C1163 a_n1500_n60543# a_n1500_n61779# 3.11f
C1164 w_n1594_n60546# a_n1500_n60543# 1.65f
C1165 w_n1594_n63018# a_n1500_n63015# 1.65f
C1166 a_n1500_3729# a_n1500_2493# 3.11f
C1167 w_n1594_46986# a_1500_47086# 0.0187f
C1168 a_n1558_n45614# a_n1558_n46850# 0.0105f
C1169 w_n1594_n13578# a_1500_n12242# 0.0023f
C1170 a_n1500_6201# w_n1594_4962# 0.0172f
C1171 a_1500_21130# a_1500_19894# 0.0105f
C1172 a_n1500_3729# w_n1594_4962# 0.0172f
C1173 a_n1558_47086# w_n1594_48222# 0.0023f
C1174 w_n1594_n34590# a_1500_n33254# 0.0023f
C1175 a_1500_32254# w_n1594_33390# 0.0023f
C1176 a_n1500_n42003# a_1500_n41906# 0.217f
C1177 a_1500_22366# w_n1594_21030# 0.0023f
C1178 w_n1594_1254# a_n1558_118# 0.0023f
C1179 w_n1594_n2454# a_n1558_n1118# 0.0023f
C1180 a_n1500_39573# a_n1558_39670# 0.217f
C1181 a_n1500_n2451# a_n1558_n2354# 0.217f
C1182 a_n1558_n53030# w_n1594_n51894# 0.0023f
C1183 a_n1500_40809# w_n1594_42042# 0.0172f
C1184 a_1500_32254# a_1500_31018# 0.0105f
C1185 w_n1594_59346# a_n1558_60682# 0.0023f
C1186 a_n1558_44614# w_n1594_45750# 0.0023f
C1187 w_n1594_37098# a_1500_38434# 0.0023f
C1188 a_n1558_2590# a_n1558_1354# 0.0105f
C1189 w_n1594_45750# a_n1500_44517# 0.0172f
C1190 a_n1500_60585# a_n1558_60682# 0.217f
C1191 a_n1500_42045# w_n1594_40806# 0.0172f
C1192 w_n1594_3726# a_n1500_4965# 0.0172f
C1193 a_n1558_50794# a_n1558_52030# 0.0105f
C1194 a_1500_50794# a_n1500_50697# 0.217f
C1195 a_n1558_n36962# w_n1594_n37062# 0.0187f
C1196 a_n1558_n23366# w_n1594_n23466# 0.0187f
C1197 a_1500_24838# a_n1500_24741# 0.217f
C1198 a_n1500_7437# w_n1594_6198# 0.0172f
C1199 a_n1500_n51891# w_n1594_n53130# 0.0172f
C1200 a_n1558_n17186# a_n1500_n17283# 0.217f
C1201 a_n1500_n33351# w_n1594_n32118# 0.0172f
C1202 a_1500_45850# a_1500_47086# 0.0105f
C1203 w_n1594_n56838# a_n1558_n56738# 0.0187f
C1204 a_1500_n32018# w_n1594_n33354# 0.0023f
C1205 w_n1594_n54366# a_n1558_n53030# 0.0023f
C1206 a_n1500_28449# w_n1594_28446# 1.65f
C1207 a_n1500_n35823# a_n1500_n37059# 3.11f
C1208 a_1500_7534# w_n1594_8670# 0.0023f
C1209 a_n1558_n44378# a_n1558_n43142# 0.0105f
C1210 w_n1594_n42006# a_n1558_n41906# 0.0187f
C1211 w_n1594_n43242# a_n1500_n42003# 0.0172f
C1212 a_1500_29782# w_n1594_28446# 0.0023f
C1213 a_n1558_n29546# w_n1594_n29646# 0.0187f
C1214 a_n1558_n4826# a_n1558_n3590# 0.0105f
C1215 a_n1558_n12242# w_n1594_n13578# 0.0023f
C1216 a_n1500_21# w_n1594_18# 1.65f
C1217 a_1500_26074# w_n1594_24738# 0.0023f
C1218 w_n1594_n61782# a_n1500_n60543# 0.0172f
C1219 w_n1594_55638# a_n1500_54405# 0.0172f
C1220 a_n1500_13617# w_n1594_13614# 1.65f
C1221 a_n1500_16089# w_n1594_17322# 0.0172f
C1222 a_1500_55738# a_1500_56974# 0.0105f
C1223 w_n1594_n58074# a_n1558_n57974# 0.0187f
C1224 a_1500_n20894# w_n1594_n20994# 0.0187f
C1225 a_n1558_n17186# w_n1594_n18522# 0.0023f
C1226 w_n1594_35862# a_1500_37198# 0.0023f
C1227 a_1500_n14714# w_n1594_n14814# 0.0187f
C1228 w_n1594_35862# a_n1558_37198# 0.0023f
C1229 a_n1500_n46947# w_n1594_n46950# 1.65f
C1230 w_n1594_n20994# a_n1558_n20894# 0.0187f
C1231 a_n1500_21033# w_n1594_21030# 1.65f
C1232 a_n1500_14853# a_n1500_16089# 3.11f
C1233 a_n1558_n39434# w_n1594_n38298# 0.0023f
C1234 a_1500_n17186# a_1500_n18422# 0.0105f
C1235 w_n1594_n63018# a_n1500_n61779# 0.0172f
C1236 a_n1500_n45711# a_1500_n45614# 0.217f
C1237 a_1500_34726# w_n1594_35862# 0.0023f
C1238 a_1500_45850# w_n1594_46986# 0.0023f
C1239 w_n1594_n29646# a_n1500_n28407# 0.0172f
C1240 a_n1500_n16047# a_n1558_n15950# 0.217f
C1241 a_n1500_n54363# a_n1558_n54266# 0.217f
C1242 a_1500_n53030# a_1500_n54266# 0.0105f
C1243 a_n1558_43378# a_n1558_44614# 0.0105f
C1244 a_n1558_18658# w_n1594_17322# 0.0023f
C1245 a_1500_n50558# a_1500_n51794# 0.0105f
C1246 a_n1558_59446# a_n1558_60682# 0.0105f
C1247 a_n1500_22269# a_n1500_23505# 3.11f
C1248 w_n1594_35862# a_n1558_34726# 0.0023f
C1249 w_n1594_n59310# a_n1558_n60446# 0.0023f
C1250 a_n1558_n40670# a_n1558_n41906# 0.0105f
C1251 a_n1500_n9867# w_n1594_n11106# 0.0172f
C1252 a_1500_n36962# w_n1594_n35826# 0.0023f
C1253 a_1500_n48086# a_1500_n49322# 0.0105f
C1254 w_n1594_n2454# a_n1558_n3590# 0.0023f
C1255 a_n1500_n49419# a_n1558_n49322# 0.217f
C1256 a_n1500_n25935# a_n1500_n24699# 3.11f
C1257 a_n1558_n8534# w_n1594_n8634# 0.0187f
C1258 a_n1558_n51794# w_n1594_n51894# 0.0187f
C1259 a_n1500_51933# w_n1594_53166# 0.0172f
C1260 w_n1594_n24702# a_1500_n25838# 0.0023f
C1261 w_n1594_4962# a_1500_6298# 0.0023f
C1262 w_n1594_13614# a_1500_14950# 0.0023f
C1263 a_1500_33490# w_n1594_32154# 0.0023f
C1264 w_n1594_n1218# a_n1558_n2354# 0.0023f
C1265 a_n1500_n3687# a_n1500_n4923# 3.11f
C1266 a_n1500_29685# w_n1594_29682# 1.65f
C1267 a_n1500_49461# w_n1594_48222# 0.0172f
C1268 w_n1594_11142# a_n1558_10006# 0.0023f
C1269 w_n1594_3726# a_1500_3826# 0.0187f
C1270 a_n1558_54502# w_n1594_53166# 0.0023f
C1271 a_n1558_13714# w_n1594_13614# 0.0187f
C1272 a_n1558_42142# w_n1594_42042# 0.0187f
C1273 w_n1594_48222# a_n1558_49558# 0.0023f
C1274 a_n1500_58113# a_n1558_58210# 0.217f
C1275 w_n1594_9906# a_n1500_8673# 0.0172f
C1276 w_n1594_4962# a_n1558_6298# 0.0023f
C1277 a_n1500_n23463# a_n1558_n23366# 0.217f
C1278 a_n1558_n35726# w_n1594_n37062# 0.0023f
C1279 w_n1594_n8634# a_n1558_n7298# 0.0023f
C1280 a_1500_53266# a_1500_54502# 0.0105f
C1281 a_n1558_n39434# a_n1558_n40670# 0.0105f
C1282 a_n1558_43378# a_n1500_43281# 0.217f
C1283 w_n1594_n9870# a_n1558_n9770# 0.0187f
C1284 a_n1500_n32115# w_n1594_n32118# 1.65f
C1285 a_n1558_47086# a_n1500_46989# 0.217f
C1286 w_n1594_n56838# a_n1558_n55502# 0.0023f
C1287 a_n1558_27310# a_n1558_26074# 0.0105f
C1288 a_n1500_16089# a_n1500_17325# 3.11f
C1289 w_n1594_58110# a_n1558_58210# 0.0187f
C1290 w_n1594_56874# a_n1558_55738# 0.0023f
C1291 a_n1500_6201# a_n1500_7437# 3.11f
C1292 a_n1558_24838# a_n1500_24741# 0.217f
C1293 a_n1558_2590# w_n1594_3726# 0.0023f
C1294 w_n1594_n42006# a_n1558_n40670# 0.0023f
C1295 a_n1500_n44475# w_n1594_n44478# 1.65f
C1296 a_n1558_33490# w_n1594_32154# 0.0023f
C1297 a_n1558_n28310# w_n1594_n29646# 0.0023f
C1298 a_n1500_7437# w_n1594_8670# 0.0172f
C1299 a_1500_7534# a_1500_6298# 0.0105f
C1300 a_n1558_n38198# a_n1558_n39434# 0.0105f
C1301 a_n1558_n17186# w_n1594_n17286# 0.0187f
C1302 w_n1594_n58074# a_n1558_n56738# 0.0023f
C1303 a_1500_23602# w_n1594_22266# 0.0023f
C1304 a_1500_48322# a_n1500_48225# 0.217f
C1305 a_n1558_n22130# a_n1500_n22227# 0.217f
C1306 a_n1500_n45711# w_n1594_n46950# 0.0172f
C1307 a_n1558_2590# a_n1558_3826# 0.0105f
C1308 a_n1500_21033# a_n1500_19797# 3.11f
C1309 a_n1500_1257# a_n1500_2493# 3.11f
C1310 a_n1558_n24602# w_n1594_n23466# 0.0023f
C1311 a_n1558_47086# a_n1558_45850# 0.0105f
C1312 a_1500_12478# a_1500_13714# 0.0105f
C1313 a_1500_2590# a_1500_3826# 0.0105f
C1314 a_1500_19894# a_1500_18658# 0.0105f
C1315 a_1500_26074# a_n1500_25977# 0.217f
C1316 a_n1500_n6159# a_n1558_n6062# 0.217f
C1317 a_n1558_n38198# w_n1594_n38298# 0.0187f
C1318 a_n1500_n7395# w_n1594_n6162# 0.0172f
C1319 a_n1558_n44378# a_n1558_n45614# 0.0105f
C1320 a_1500_55738# a_n1500_55641# 0.217f
C1321 a_n1558_45850# w_n1594_44514# 0.0023f
C1322 a_n1558_n49322# w_n1594_n48186# 0.0023f
C1323 a_n1500_n20991# w_n1594_n20994# 1.65f
C1324 a_1500_n4826# w_n1594_n3690# 0.0023f
C1325 a_1500_118# a_1500_1354# 0.0105f
C1326 a_n1500_n63015# a_1500_n62918# 0.217f
C1327 a_n1500_n40767# a_1500_n40670# 0.217f
C1328 w_n1594_n59310# a_n1558_n59210# 0.0187f
C1329 a_n1500_24741# a_n1500_23505# 3.11f
C1330 a_1500_7534# a_1500_8770# 0.0105f
C1331 a_1500_n35726# w_n1594_n35826# 0.0187f
C1332 w_n1594_48222# a_n1500_48225# 1.65f
C1333 a_n1500_n33351# a_n1500_n34587# 3.11f
C1334 a_n1558_39670# w_n1594_40806# 0.0023f
C1335 w_n1594_n14814# a_1500_n15950# 0.0023f
C1336 a_n1558_50794# a_n1558_49558# 0.0105f
C1337 a_1500_5062# a_1500_6298# 0.0105f
C1338 a_n1500_24741# w_n1594_24738# 1.65f
C1339 a_n1558_n11006# a_n1558_n9770# 0.0105f
C1340 a_n1558_27310# a_n1558_28546# 0.0105f
C1341 a_n1558_n50558# w_n1594_n49422# 0.0023f
C1342 w_n1594_55638# a_1500_54502# 0.0023f
C1343 a_n1500_n56835# a_n1500_n58071# 3.11f
C1344 a_n1500_n50655# w_n1594_n50658# 1.65f
C1345 a_n1500_1257# a_1500_1354# 0.217f
C1346 a_1500_n2354# a_n1500_n2451# 0.217f
C1347 a_1500_40906# w_n1594_42042# 0.0023f
C1348 w_n1594_n30882# a_n1500_n30879# 1.65f
C1349 a_n1500_n13575# a_n1500_n12339# 3.11f
C1350 a_n1558_5062# a_n1500_4965# 0.217f
C1351 w_n1594_n3690# a_n1558_n3590# 0.0187f
C1352 a_n1500_n39531# a_1500_n39434# 0.217f
C1353 w_n1594_61818# a_n1558_60682# 0.0023f
C1354 w_n1594_54402# a_n1558_53266# 0.0023f
C1355 a_n1500_51933# w_n1594_51930# 1.65f
C1356 a_1500_n3590# w_n1594_n2454# 0.0023f
C1357 a_1500_19894# w_n1594_21030# 0.0023f
C1358 w_n1594_n55602# a_1500_n56738# 0.0023f
C1359 a_1500_26074# w_n1594_27210# 0.0023f
C1360 a_n1558_32254# a_n1558_31018# 0.0105f
C1361 a_n1558_32254# a_n1500_32157# 0.217f
C1362 a_n1500_n59307# a_n1558_n59210# 0.217f
C1363 a_1500_49558# a_1500_48322# 0.0105f
C1364 a_n1500_45753# w_n1594_45750# 1.65f
C1365 a_n1500_n43239# w_n1594_n44478# 0.0172f
C1366 a_1500_16186# w_n1594_16086# 0.0187f
C1367 a_n1500_21# w_n1594_n1218# 0.0172f
C1368 a_n1558_54502# a_n1558_53266# 0.0105f
C1369 a_1500_21130# w_n1594_21030# 0.0187f
C1370 a_n1500_58113# a_1500_58210# 0.217f
C1371 a_1500_53266# a_n1500_53169# 0.217f
C1372 a_n1500_29685# a_n1558_29782# 0.217f
C1373 a_n1500_n38295# a_1500_n38198# 0.217f
C1374 a_1500_14950# w_n1594_16086# 0.0023f
C1375 a_n1500_3729# w_n1594_2490# 0.0172f
C1376 a_n1500_35865# w_n1594_34626# 0.0172f
C1377 a_n1500_n29643# a_n1500_n30879# 3.11f
C1378 a_n1500_39573# a_1500_39670# 0.217f
C1379 w_n1594_58110# a_1500_58210# 0.0187f
C1380 w_n1594_56874# a_n1500_58113# 0.0172f
C1381 w_n1594_54402# a_n1500_54405# 1.65f
C1382 a_n1558_n46850# w_n1594_n45714# 0.0023f
C1383 w_n1594_60582# a_n1500_59349# 0.0172f
C1384 a_n1500_n3687# a_n1500_n2451# 3.11f
C1385 w_n1594_n34590# a_n1500_n35823# 0.0172f
C1386 a_n1558_n36962# w_n1594_n38298# 0.0023f
C1387 a_n1558_n13478# a_n1558_n14714# 0.0105f
C1388 a_n1558_27310# w_n1594_27210# 0.0187f
C1389 a_1500_49558# w_n1594_48222# 0.0023f
C1390 a_1500_n34490# a_1500_n35726# 0.0105f
C1391 a_n1558_54502# a_n1500_54405# 0.217f
C1392 a_n1558_n25838# w_n1594_n27174# 0.0023f
C1393 a_n1558_19894# a_n1558_21130# 0.0105f
C1394 a_n1558_n48086# w_n1594_n48186# 0.0187f
C1395 a_1500_33490# w_n1594_34626# 0.0023f
C1396 a_n1500_n53127# a_n1558_n53030# 0.217f
C1397 a_1500_n51794# a_1500_n53030# 0.0105f
C1398 a_n1558_n61682# a_n1558_n62918# 0.0105f
C1399 a_n1500_37101# w_n1594_38334# 0.0172f
C1400 a_n1500_n48183# a_n1558_n48086# 0.217f
C1401 w_n1594_n20994# a_n1558_n19658# 0.0023f
C1402 a_1500_n46850# a_1500_n48086# 0.0105f
C1403 w_n1594_45750# a_1500_47086# 0.0023f
C1404 a_n1558_11242# a_n1558_10006# 0.0105f
C1405 a_1500_13714# w_n1594_14850# 0.0023f
C1406 a_n1558_16186# w_n1594_14850# 0.0023f
C1407 a_n1500_n7395# a_n1558_n7298# 0.217f
C1408 a_n1500_21# a_n1500_n1215# 3.11f
C1409 a_n1558_n49322# w_n1594_n49422# 0.0187f
C1410 w_n1594_60582# a_1500_59446# 0.0023f
C1411 w_n1594_60582# a_1500_60682# 0.0187f
C1412 a_1500_n2354# a_1500_n1118# 0.0105f
C1413 w_n1594_48222# a_n1558_48322# 0.0187f
C1414 a_n1500_n49419# w_n1594_n50658# 0.0172f
C1415 a_n1500_21033# w_n1594_19794# 0.0172f
C1416 a_1500_52030# a_1500_53266# 0.0105f
C1417 a_1500_42142# a_1500_43378# 0.0105f
C1418 w_n1594_n18522# a_n1558_n19658# 0.0023f
C1419 a_1500_n62918# VSUBS 0.638f
C1420 a_n1558_n62918# VSUBS 0.638f
C1421 a_n1500_n63015# VSUBS 5.03f
C1422 a_1500_n61682# VSUBS 0.625f
C1423 a_n1558_n61682# VSUBS 0.625f
C1424 a_n1500_n61779# VSUBS 3.31f
C1425 a_1500_n60446# VSUBS 0.625f
C1426 a_n1558_n60446# VSUBS 0.625f
C1427 a_n1500_n60543# VSUBS 3.31f
C1428 a_1500_n59210# VSUBS 0.625f
C1429 a_n1558_n59210# VSUBS 0.625f
C1430 a_n1500_n59307# VSUBS 3.31f
C1431 a_1500_n57974# VSUBS 0.625f
C1432 a_n1558_n57974# VSUBS 0.625f
C1433 a_n1500_n58071# VSUBS 3.31f
C1434 a_1500_n56738# VSUBS 0.625f
C1435 a_n1558_n56738# VSUBS 0.625f
C1436 a_n1500_n56835# VSUBS 3.31f
C1437 a_1500_n55502# VSUBS 0.625f
C1438 a_n1558_n55502# VSUBS 0.625f
C1439 a_n1500_n55599# VSUBS 3.31f
C1440 a_1500_n54266# VSUBS 0.625f
C1441 a_n1558_n54266# VSUBS 0.625f
C1442 a_n1500_n54363# VSUBS 3.31f
C1443 a_1500_n53030# VSUBS 0.625f
C1444 a_n1558_n53030# VSUBS 0.625f
C1445 a_n1500_n53127# VSUBS 3.31f
C1446 a_1500_n51794# VSUBS 0.625f
C1447 a_n1558_n51794# VSUBS 0.625f
C1448 a_n1500_n51891# VSUBS 3.31f
C1449 a_1500_n50558# VSUBS 0.625f
C1450 a_n1558_n50558# VSUBS 0.625f
C1451 a_n1500_n50655# VSUBS 3.31f
C1452 a_1500_n49322# VSUBS 0.625f
C1453 a_n1558_n49322# VSUBS 0.625f
C1454 a_n1500_n49419# VSUBS 3.31f
C1455 a_1500_n48086# VSUBS 0.625f
C1456 a_n1558_n48086# VSUBS 0.625f
C1457 a_n1500_n48183# VSUBS 3.31f
C1458 a_1500_n46850# VSUBS 0.625f
C1459 a_n1558_n46850# VSUBS 0.625f
C1460 a_n1500_n46947# VSUBS 3.31f
C1461 a_1500_n45614# VSUBS 0.625f
C1462 a_n1558_n45614# VSUBS 0.625f
C1463 a_n1500_n45711# VSUBS 3.31f
C1464 a_1500_n44378# VSUBS 0.625f
C1465 a_n1558_n44378# VSUBS 0.625f
C1466 a_n1500_n44475# VSUBS 3.31f
C1467 a_1500_n43142# VSUBS 0.625f
C1468 a_n1558_n43142# VSUBS 0.625f
C1469 a_n1500_n43239# VSUBS 3.31f
C1470 a_1500_n41906# VSUBS 0.625f
C1471 a_n1558_n41906# VSUBS 0.625f
C1472 a_n1500_n42003# VSUBS 3.31f
C1473 a_1500_n40670# VSUBS 0.625f
C1474 a_n1558_n40670# VSUBS 0.625f
C1475 a_n1500_n40767# VSUBS 3.31f
C1476 a_1500_n39434# VSUBS 0.625f
C1477 a_n1558_n39434# VSUBS 0.625f
C1478 a_n1500_n39531# VSUBS 3.31f
C1479 a_1500_n38198# VSUBS 0.625f
C1480 a_n1558_n38198# VSUBS 0.625f
C1481 a_n1500_n38295# VSUBS 3.31f
C1482 a_1500_n36962# VSUBS 0.625f
C1483 a_n1558_n36962# VSUBS 0.625f
C1484 a_n1500_n37059# VSUBS 3.31f
C1485 a_1500_n35726# VSUBS 0.625f
C1486 a_n1558_n35726# VSUBS 0.625f
C1487 a_n1500_n35823# VSUBS 3.31f
C1488 a_1500_n34490# VSUBS 0.625f
C1489 a_n1558_n34490# VSUBS 0.625f
C1490 a_n1500_n34587# VSUBS 3.31f
C1491 a_1500_n33254# VSUBS 0.625f
C1492 a_n1558_n33254# VSUBS 0.625f
C1493 a_n1500_n33351# VSUBS 3.31f
C1494 a_1500_n32018# VSUBS 0.625f
C1495 a_n1558_n32018# VSUBS 0.625f
C1496 a_n1500_n32115# VSUBS 3.31f
C1497 a_1500_n30782# VSUBS 0.625f
C1498 a_n1558_n30782# VSUBS 0.625f
C1499 a_n1500_n30879# VSUBS 3.31f
C1500 a_1500_n29546# VSUBS 0.625f
C1501 a_n1558_n29546# VSUBS 0.625f
C1502 a_n1500_n29643# VSUBS 3.31f
C1503 a_1500_n28310# VSUBS 0.625f
C1504 a_n1558_n28310# VSUBS 0.625f
C1505 a_n1500_n28407# VSUBS 3.31f
C1506 a_1500_n27074# VSUBS 0.625f
C1507 a_n1558_n27074# VSUBS 0.625f
C1508 a_n1500_n27171# VSUBS 3.31f
C1509 a_1500_n25838# VSUBS 0.625f
C1510 a_n1558_n25838# VSUBS 0.625f
C1511 a_n1500_n25935# VSUBS 3.31f
C1512 a_1500_n24602# VSUBS 0.625f
C1513 a_n1558_n24602# VSUBS 0.625f
C1514 a_n1500_n24699# VSUBS 3.31f
C1515 a_1500_n23366# VSUBS 0.625f
C1516 a_n1558_n23366# VSUBS 0.625f
C1517 a_n1500_n23463# VSUBS 3.31f
C1518 a_1500_n22130# VSUBS 0.625f
C1519 a_n1558_n22130# VSUBS 0.625f
C1520 a_n1500_n22227# VSUBS 3.31f
C1521 a_1500_n20894# VSUBS 0.625f
C1522 a_n1558_n20894# VSUBS 0.625f
C1523 a_n1500_n20991# VSUBS 3.31f
C1524 a_1500_n19658# VSUBS 0.625f
C1525 a_n1558_n19658# VSUBS 0.625f
C1526 a_n1500_n19755# VSUBS 3.31f
C1527 a_1500_n18422# VSUBS 0.625f
C1528 a_n1558_n18422# VSUBS 0.625f
C1529 a_n1500_n18519# VSUBS 3.31f
C1530 a_1500_n17186# VSUBS 0.625f
C1531 a_n1558_n17186# VSUBS 0.625f
C1532 a_n1500_n17283# VSUBS 3.31f
C1533 a_1500_n15950# VSUBS 0.625f
C1534 a_n1558_n15950# VSUBS 0.625f
C1535 a_n1500_n16047# VSUBS 3.31f
C1536 a_1500_n14714# VSUBS 0.625f
C1537 a_n1558_n14714# VSUBS 0.625f
C1538 a_n1500_n14811# VSUBS 3.31f
C1539 a_1500_n13478# VSUBS 0.625f
C1540 a_n1558_n13478# VSUBS 0.625f
C1541 a_n1500_n13575# VSUBS 3.31f
C1542 a_1500_n12242# VSUBS 0.625f
C1543 a_n1558_n12242# VSUBS 0.625f
C1544 a_n1500_n12339# VSUBS 3.31f
C1545 a_1500_n11006# VSUBS 0.625f
C1546 a_n1558_n11006# VSUBS 0.625f
C1547 a_n1500_n11103# VSUBS 3.31f
C1548 a_1500_n9770# VSUBS 0.625f
C1549 a_n1558_n9770# VSUBS 0.625f
C1550 a_n1500_n9867# VSUBS 3.31f
C1551 a_1500_n8534# VSUBS 0.625f
C1552 a_n1558_n8534# VSUBS 0.625f
C1553 a_n1500_n8631# VSUBS 3.31f
C1554 a_1500_n7298# VSUBS 0.625f
C1555 a_n1558_n7298# VSUBS 0.625f
C1556 a_n1500_n7395# VSUBS 3.31f
C1557 a_1500_n6062# VSUBS 0.625f
C1558 a_n1558_n6062# VSUBS 0.625f
C1559 a_n1500_n6159# VSUBS 3.31f
C1560 a_1500_n4826# VSUBS 0.625f
C1561 a_n1558_n4826# VSUBS 0.625f
C1562 a_n1500_n4923# VSUBS 3.31f
C1563 a_1500_n3590# VSUBS 0.625f
C1564 a_n1558_n3590# VSUBS 0.625f
C1565 a_n1500_n3687# VSUBS 3.31f
C1566 a_1500_n2354# VSUBS 0.625f
C1567 a_n1558_n2354# VSUBS 0.625f
C1568 a_n1500_n2451# VSUBS 3.31f
C1569 a_1500_n1118# VSUBS 0.625f
C1570 a_n1558_n1118# VSUBS 0.625f
C1571 a_n1500_n1215# VSUBS 3.31f
C1572 a_1500_118# VSUBS 0.625f
C1573 a_n1558_118# VSUBS 0.625f
C1574 a_n1500_21# VSUBS 3.31f
C1575 a_1500_1354# VSUBS 0.625f
C1576 a_n1558_1354# VSUBS 0.625f
C1577 a_n1500_1257# VSUBS 3.31f
C1578 a_1500_2590# VSUBS 0.625f
C1579 a_n1558_2590# VSUBS 0.625f
C1580 a_n1500_2493# VSUBS 3.31f
C1581 a_1500_3826# VSUBS 0.625f
C1582 a_n1558_3826# VSUBS 0.625f
C1583 a_n1500_3729# VSUBS 3.31f
C1584 a_1500_5062# VSUBS 0.625f
C1585 a_n1558_5062# VSUBS 0.625f
C1586 a_n1500_4965# VSUBS 3.31f
C1587 a_1500_6298# VSUBS 0.625f
C1588 a_n1558_6298# VSUBS 0.625f
C1589 a_n1500_6201# VSUBS 3.31f
C1590 a_1500_7534# VSUBS 0.625f
C1591 a_n1558_7534# VSUBS 0.625f
C1592 a_n1500_7437# VSUBS 3.31f
C1593 a_1500_8770# VSUBS 0.625f
C1594 a_n1558_8770# VSUBS 0.625f
C1595 a_n1500_8673# VSUBS 3.31f
C1596 a_1500_10006# VSUBS 0.625f
C1597 a_n1558_10006# VSUBS 0.625f
C1598 a_n1500_9909# VSUBS 3.31f
C1599 a_1500_11242# VSUBS 0.625f
C1600 a_n1558_11242# VSUBS 0.625f
C1601 a_n1500_11145# VSUBS 3.31f
C1602 a_1500_12478# VSUBS 0.625f
C1603 a_n1558_12478# VSUBS 0.625f
C1604 a_n1500_12381# VSUBS 3.31f
C1605 a_1500_13714# VSUBS 0.625f
C1606 a_n1558_13714# VSUBS 0.625f
C1607 a_n1500_13617# VSUBS 3.31f
C1608 a_1500_14950# VSUBS 0.625f
C1609 a_n1558_14950# VSUBS 0.625f
C1610 a_n1500_14853# VSUBS 3.31f
C1611 a_1500_16186# VSUBS 0.625f
C1612 a_n1558_16186# VSUBS 0.625f
C1613 a_n1500_16089# VSUBS 3.31f
C1614 a_1500_17422# VSUBS 0.625f
C1615 a_n1558_17422# VSUBS 0.625f
C1616 a_n1500_17325# VSUBS 3.31f
C1617 a_1500_18658# VSUBS 0.625f
C1618 a_n1558_18658# VSUBS 0.625f
C1619 a_n1500_18561# VSUBS 3.31f
C1620 a_1500_19894# VSUBS 0.625f
C1621 a_n1558_19894# VSUBS 0.625f
C1622 a_n1500_19797# VSUBS 3.31f
C1623 a_1500_21130# VSUBS 0.625f
C1624 a_n1558_21130# VSUBS 0.625f
C1625 a_n1500_21033# VSUBS 3.31f
C1626 a_1500_22366# VSUBS 0.625f
C1627 a_n1558_22366# VSUBS 0.625f
C1628 a_n1500_22269# VSUBS 3.31f
C1629 a_1500_23602# VSUBS 0.625f
C1630 a_n1558_23602# VSUBS 0.625f
C1631 a_n1500_23505# VSUBS 3.31f
C1632 a_1500_24838# VSUBS 0.625f
C1633 a_n1558_24838# VSUBS 0.625f
C1634 a_n1500_24741# VSUBS 3.31f
C1635 a_1500_26074# VSUBS 0.625f
C1636 a_n1558_26074# VSUBS 0.625f
C1637 a_n1500_25977# VSUBS 3.31f
C1638 a_1500_27310# VSUBS 0.625f
C1639 a_n1558_27310# VSUBS 0.625f
C1640 a_n1500_27213# VSUBS 3.31f
C1641 a_1500_28546# VSUBS 0.625f
C1642 a_n1558_28546# VSUBS 0.625f
C1643 a_n1500_28449# VSUBS 3.31f
C1644 a_1500_29782# VSUBS 0.625f
C1645 a_n1558_29782# VSUBS 0.625f
C1646 a_n1500_29685# VSUBS 3.31f
C1647 a_1500_31018# VSUBS 0.625f
C1648 a_n1558_31018# VSUBS 0.625f
C1649 a_n1500_30921# VSUBS 3.31f
C1650 a_1500_32254# VSUBS 0.625f
C1651 a_n1558_32254# VSUBS 0.625f
C1652 a_n1500_32157# VSUBS 3.31f
C1653 a_1500_33490# VSUBS 0.625f
C1654 a_n1558_33490# VSUBS 0.625f
C1655 a_n1500_33393# VSUBS 3.31f
C1656 a_1500_34726# VSUBS 0.625f
C1657 a_n1558_34726# VSUBS 0.625f
C1658 a_n1500_34629# VSUBS 3.31f
C1659 a_1500_35962# VSUBS 0.625f
C1660 a_n1558_35962# VSUBS 0.625f
C1661 a_n1500_35865# VSUBS 3.31f
C1662 a_1500_37198# VSUBS 0.625f
C1663 a_n1558_37198# VSUBS 0.625f
C1664 a_n1500_37101# VSUBS 3.31f
C1665 a_1500_38434# VSUBS 0.625f
C1666 a_n1558_38434# VSUBS 0.625f
C1667 a_n1500_38337# VSUBS 3.31f
C1668 a_1500_39670# VSUBS 0.625f
C1669 a_n1558_39670# VSUBS 0.625f
C1670 a_n1500_39573# VSUBS 3.31f
C1671 a_1500_40906# VSUBS 0.625f
C1672 a_n1558_40906# VSUBS 0.625f
C1673 a_n1500_40809# VSUBS 3.31f
C1674 a_1500_42142# VSUBS 0.625f
C1675 a_n1558_42142# VSUBS 0.625f
C1676 a_n1500_42045# VSUBS 3.31f
C1677 a_1500_43378# VSUBS 0.625f
C1678 a_n1558_43378# VSUBS 0.625f
C1679 a_n1500_43281# VSUBS 3.31f
C1680 a_1500_44614# VSUBS 0.625f
C1681 a_n1558_44614# VSUBS 0.625f
C1682 a_n1500_44517# VSUBS 3.31f
C1683 a_1500_45850# VSUBS 0.625f
C1684 a_n1558_45850# VSUBS 0.625f
C1685 a_n1500_45753# VSUBS 3.31f
C1686 a_1500_47086# VSUBS 0.625f
C1687 a_n1558_47086# VSUBS 0.625f
C1688 a_n1500_46989# VSUBS 3.31f
C1689 a_1500_48322# VSUBS 0.625f
C1690 a_n1558_48322# VSUBS 0.625f
C1691 a_n1500_48225# VSUBS 3.31f
C1692 a_1500_49558# VSUBS 0.625f
C1693 a_n1558_49558# VSUBS 0.625f
C1694 a_n1500_49461# VSUBS 3.31f
C1695 a_1500_50794# VSUBS 0.625f
C1696 a_n1558_50794# VSUBS 0.625f
C1697 a_n1500_50697# VSUBS 3.31f
C1698 a_1500_52030# VSUBS 0.625f
C1699 a_n1558_52030# VSUBS 0.625f
C1700 a_n1500_51933# VSUBS 3.31f
C1701 a_1500_53266# VSUBS 0.625f
C1702 a_n1558_53266# VSUBS 0.625f
C1703 a_n1500_53169# VSUBS 3.31f
C1704 a_1500_54502# VSUBS 0.625f
C1705 a_n1558_54502# VSUBS 0.625f
C1706 a_n1500_54405# VSUBS 3.31f
C1707 a_1500_55738# VSUBS 0.625f
C1708 a_n1558_55738# VSUBS 0.625f
C1709 a_n1500_55641# VSUBS 3.31f
C1710 a_1500_56974# VSUBS 0.625f
C1711 a_n1558_56974# VSUBS 0.625f
C1712 a_n1500_56877# VSUBS 3.31f
C1713 a_1500_58210# VSUBS 0.625f
C1714 a_n1558_58210# VSUBS 0.625f
C1715 a_n1500_58113# VSUBS 3.31f
C1716 a_1500_59446# VSUBS 0.625f
C1717 a_n1558_59446# VSUBS 0.625f
C1718 a_n1500_59349# VSUBS 3.31f
C1719 a_1500_60682# VSUBS 0.625f
C1720 a_n1558_60682# VSUBS 0.625f
C1721 a_n1500_60585# VSUBS 3.31f
C1722 a_1500_61918# VSUBS 0.638f
C1723 a_n1558_61918# VSUBS 0.638f
C1724 a_n1500_61821# VSUBS 5.03f
C1725 w_n1594_n63018# VSUBS 11.5f
C1726 w_n1594_n61782# VSUBS 11.5f
C1727 w_n1594_n60546# VSUBS 11.5f
C1728 w_n1594_n59310# VSUBS 11.5f
C1729 w_n1594_n58074# VSUBS 11.5f
C1730 w_n1594_n56838# VSUBS 11.5f
C1731 w_n1594_n55602# VSUBS 11.5f
C1732 w_n1594_n54366# VSUBS 11.5f
C1733 w_n1594_n53130# VSUBS 11.5f
C1734 w_n1594_n51894# VSUBS 11.5f
C1735 w_n1594_n50658# VSUBS 11.5f
C1736 w_n1594_n49422# VSUBS 11.5f
C1737 w_n1594_n48186# VSUBS 11.5f
C1738 w_n1594_n46950# VSUBS 11.5f
C1739 w_n1594_n45714# VSUBS 11.5f
C1740 w_n1594_n44478# VSUBS 11.5f
C1741 w_n1594_n43242# VSUBS 11.5f
C1742 w_n1594_n42006# VSUBS 11.5f
C1743 w_n1594_n40770# VSUBS 11.5f
C1744 w_n1594_n39534# VSUBS 11.5f
C1745 w_n1594_n38298# VSUBS 11.5f
C1746 w_n1594_n37062# VSUBS 11.5f
C1747 w_n1594_n35826# VSUBS 11.5f
C1748 w_n1594_n34590# VSUBS 11.5f
C1749 w_n1594_n33354# VSUBS 11.5f
C1750 w_n1594_n32118# VSUBS 11.5f
C1751 w_n1594_n30882# VSUBS 11.5f
C1752 w_n1594_n29646# VSUBS 11.5f
C1753 w_n1594_n28410# VSUBS 11.5f
C1754 w_n1594_n27174# VSUBS 11.5f
C1755 w_n1594_n25938# VSUBS 11.5f
C1756 w_n1594_n24702# VSUBS 11.5f
C1757 w_n1594_n23466# VSUBS 11.5f
C1758 w_n1594_n22230# VSUBS 11.5f
C1759 w_n1594_n20994# VSUBS 11.5f
C1760 w_n1594_n19758# VSUBS 11.5f
C1761 w_n1594_n18522# VSUBS 11.5f
C1762 w_n1594_n17286# VSUBS 11.5f
C1763 w_n1594_n16050# VSUBS 11.5f
C1764 w_n1594_n14814# VSUBS 11.5f
C1765 w_n1594_n13578# VSUBS 11.5f
C1766 w_n1594_n12342# VSUBS 11.5f
C1767 w_n1594_n11106# VSUBS 11.5f
C1768 w_n1594_n9870# VSUBS 11.5f
C1769 w_n1594_n8634# VSUBS 11.5f
C1770 w_n1594_n7398# VSUBS 11.5f
C1771 w_n1594_n6162# VSUBS 11.5f
C1772 w_n1594_n4926# VSUBS 11.5f
C1773 w_n1594_n3690# VSUBS 11.5f
C1774 w_n1594_n2454# VSUBS 11.5f
C1775 w_n1594_n1218# VSUBS 11.5f
C1776 w_n1594_18# VSUBS 11.5f
C1777 w_n1594_1254# VSUBS 11.5f
C1778 w_n1594_2490# VSUBS 11.5f
C1779 w_n1594_3726# VSUBS 11.5f
C1780 w_n1594_4962# VSUBS 11.5f
C1781 w_n1594_6198# VSUBS 11.5f
C1782 w_n1594_7434# VSUBS 11.5f
C1783 w_n1594_8670# VSUBS 11.5f
C1784 w_n1594_9906# VSUBS 11.5f
C1785 w_n1594_11142# VSUBS 11.5f
C1786 w_n1594_12378# VSUBS 11.5f
C1787 w_n1594_13614# VSUBS 11.5f
C1788 w_n1594_14850# VSUBS 11.5f
C1789 w_n1594_16086# VSUBS 11.5f
C1790 w_n1594_17322# VSUBS 11.5f
C1791 w_n1594_18558# VSUBS 11.5f
C1792 w_n1594_19794# VSUBS 11.5f
C1793 w_n1594_21030# VSUBS 11.5f
C1794 w_n1594_22266# VSUBS 11.5f
C1795 w_n1594_23502# VSUBS 11.5f
C1796 w_n1594_24738# VSUBS 11.5f
C1797 w_n1594_25974# VSUBS 11.5f
C1798 w_n1594_27210# VSUBS 11.5f
C1799 w_n1594_28446# VSUBS 11.5f
C1800 w_n1594_29682# VSUBS 11.5f
C1801 w_n1594_30918# VSUBS 11.5f
C1802 w_n1594_32154# VSUBS 11.5f
C1803 w_n1594_33390# VSUBS 11.5f
C1804 w_n1594_34626# VSUBS 11.5f
C1805 w_n1594_35862# VSUBS 11.5f
C1806 w_n1594_37098# VSUBS 11.5f
C1807 w_n1594_38334# VSUBS 11.5f
C1808 w_n1594_39570# VSUBS 11.5f
C1809 w_n1594_40806# VSUBS 11.5f
C1810 w_n1594_42042# VSUBS 11.5f
C1811 w_n1594_43278# VSUBS 11.5f
C1812 w_n1594_44514# VSUBS 11.5f
C1813 w_n1594_45750# VSUBS 11.5f
C1814 w_n1594_46986# VSUBS 11.5f
C1815 w_n1594_48222# VSUBS 11.5f
C1816 w_n1594_49458# VSUBS 11.5f
C1817 w_n1594_50694# VSUBS 11.5f
C1818 w_n1594_51930# VSUBS 11.5f
C1819 w_n1594_53166# VSUBS 11.5f
C1820 w_n1594_54402# VSUBS 11.5f
C1821 w_n1594_55638# VSUBS 11.5f
C1822 w_n1594_56874# VSUBS 11.5f
C1823 w_n1594_58110# VSUBS 11.5f
C1824 w_n1594_59346# VSUBS 11.5f
C1825 w_n1594_60582# VSUBS 11.5f
C1826 w_n1594_61818# VSUBS 11.5f
.ends

.subckt sky130_fd_pr__pfet_01v8_UDMRD5 a_n558_n10388# a_n558_n7916# a_n500_5583# a_n500_n10485#
+ a_500_1972# a_n558_8152# a_n500_8055# a_500_4444# w_n594_3108# w_n594_6816# a_500_n2972#
+ a_500_736# a_500_n5444# a_n500_n597# w_n594_636# a_500_n500# a_500_9388# w_n594_n3072#
+ a_n558_1972# w_n594_n6780# w_n594_n600# a_n500_1875# a_n558_4444# w_n594_n9252#
+ a_n500_4347# a_n558_n6680# w_n594_n10488# a_n558_n9152# a_n500_n5541# a_n500_639#
+ a_500_3208# a_n500_n8013# a_500_6916# a_500_n1736# a_n558_n500# a_n558_9388# a_500_n4208#
+ w_n594_5580# a_500_n7916# w_n594_8052# w_n594_n5544# a_n558_736# a_n558_3208# w_n594_n8016#
+ a_n558_n2972# a_n558_6916# a_n558_n5444# a_n500_n1833# a_n500_6819# a_n500_n4305#
+ w_n594_1872# a_500_5680# a_n500_9291# a_n500_n3069# w_n594_4344# a_n500_n6777# a_500_8152#
+ w_n594_n1836# a_n500_n9249# a_500_n6680# w_n594_n4308# a_500_n10388# a_n500_3111#
+ a_500_n9152# a_n558_n1736# w_n594_9288# a_n558_n4208# a_n558_5680# VSUBS
X0 a_500_1972# a_n500_1875# a_n558_1972# w_n594_1872# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X1 a_500_6916# a_n500_6819# a_n558_6916# w_n594_6816# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X2 a_500_4444# a_n500_4347# a_n558_4444# w_n594_4344# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X3 a_500_n9152# a_n500_n9249# a_n558_n9152# w_n594_n9252# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X4 a_500_3208# a_n500_3111# a_n558_3208# w_n594_3108# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X5 a_500_n2972# a_n500_n3069# a_n558_n2972# w_n594_n3072# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X6 a_500_n7916# a_n500_n8013# a_n558_n7916# w_n594_n8016# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X7 a_500_9388# a_n500_9291# a_n558_9388# w_n594_9288# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X8 a_500_n5444# a_n500_n5541# a_n558_n5444# w_n594_n5544# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X9 a_500_n500# a_n500_n597# a_n558_n500# w_n594_n600# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X10 a_500_n1736# a_n500_n1833# a_n558_n1736# w_n594_n1836# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X11 a_500_n4208# a_n500_n4305# a_n558_n4208# w_n594_n4308# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X12 a_500_n10388# a_n500_n10485# a_n558_n10388# w_n594_n10488# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X13 a_500_736# a_n500_639# a_n558_736# w_n594_636# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X14 a_500_n6680# a_n500_n6777# a_n558_n6680# w_n594_n6780# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X15 a_500_5680# a_n500_5583# a_n558_5680# w_n594_5580# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X16 a_500_8152# a_n500_8055# a_n558_8152# w_n594_8052# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
C0 a_n500_n8013# a_n500_n6777# 1.03f
C1 a_n558_1972# w_n594_3108# 0.0023f
C2 a_n500_1875# a_n500_3111# 1.03f
C3 w_n594_8052# a_n500_6819# 0.00575f
C4 w_n594_n8016# a_n558_n6680# 0.0023f
C5 w_n594_n6780# a_n500_n6777# 0.593f
C6 w_n594_636# a_n558_736# 0.0187f
C7 w_n594_5580# a_n558_6916# 0.0023f
C8 a_500_n1736# a_500_n2972# 0.0105f
C9 w_n594_9288# a_n500_8055# 0.00575f
C10 a_n500_4347# a_500_4444# 0.204f
C11 w_n594_n5544# a_500_n6680# 0.0023f
C12 w_n594_636# a_500_1972# 0.0023f
C13 a_n558_n4208# a_n558_n2972# 0.0105f
C14 w_n594_9288# a_500_9388# 0.0187f
C15 a_n500_4347# w_n594_3108# 0.00575f
C16 a_500_n10388# a_n500_n10485# 0.204f
C17 a_500_5680# a_n500_5583# 0.204f
C18 a_500_6916# a_500_8152# 0.0105f
C19 w_n594_n4308# a_n500_n3069# 0.00575f
C20 a_n500_n3069# a_500_n2972# 0.204f
C21 w_n594_1872# a_n500_3111# 0.00575f
C22 a_500_n9152# a_n558_n9152# 0.0663f
C23 a_500_736# a_n558_736# 0.0663f
C24 w_n594_636# a_n558_1972# 0.0023f
C25 a_n500_5583# w_n594_6816# 0.00575f
C26 a_500_6916# a_n500_6819# 0.204f
C27 a_n558_3208# w_n594_4344# 0.0023f
C28 a_n558_n1736# w_n594_n1836# 0.0187f
C29 a_500_736# a_500_1972# 0.0105f
C30 a_500_n10388# w_n594_n10488# 0.0187f
C31 a_n500_8055# a_n558_8152# 0.204f
C32 w_n594_9288# a_n558_9388# 0.0187f
C33 w_n594_6816# a_n558_8152# 0.0023f
C34 a_500_6916# w_n594_8052# 0.0023f
C35 w_n594_n3072# a_n500_n1833# 0.00575f
C36 a_500_3208# w_n594_4344# 0.0023f
C37 a_n500_n10485# w_n594_n10488# 0.593f
C38 a_n558_n500# w_n594_n600# 0.0187f
C39 w_n594_4344# a_n558_5680# 0.0023f
C40 a_n558_6916# a_n558_8152# 0.0105f
C41 a_n500_n1833# w_n594_n600# 0.00575f
C42 a_n558_n4208# a_n558_n5444# 0.0105f
C43 w_n594_n8016# a_500_n9152# 0.0023f
C44 w_n594_n1836# a_500_n2972# 0.0023f
C45 a_n558_9388# a_n558_8152# 0.0105f
C46 w_n594_n5544# a_n500_n5541# 0.593f
C47 a_500_n10388# a_500_n9152# 0.0105f
C48 a_500_n500# a_500_n1736# 0.0105f
C49 a_n558_n7916# w_n594_n9252# 0.0023f
C50 w_n594_n3072# a_n558_n4208# 0.0023f
C51 w_n594_n5544# a_n558_n6680# 0.0023f
C52 a_n500_9291# w_n594_9288# 0.593f
C53 w_n594_n9252# a_n558_n9152# 0.0187f
C54 w_n594_3108# a_500_4444# 0.0023f
C55 a_n500_n597# a_n558_n500# 0.204f
C56 a_n558_4444# w_n594_4344# 0.0187f
C57 w_n594_n3072# a_500_n4208# 0.0023f
C58 w_n594_n4308# a_n500_n4305# 0.593f
C59 a_n500_n597# a_n500_n1833# 1.03f
C60 a_n558_n1736# a_n558_n2972# 0.0105f
C61 a_500_5680# a_500_4444# 0.0105f
C62 a_500_3208# a_n558_3208# 0.0663f
C63 a_n500_4347# a_n500_3111# 1.03f
C64 a_n500_n597# w_n594_n600# 0.593f
C65 w_n594_n10488# a_500_n9152# 0.0023f
C66 a_n558_n9152# a_n500_n9249# 0.204f
C67 w_n594_n1836# a_500_n1736# 0.0187f
C68 a_n500_n4305# a_n500_n5541# 1.03f
C69 w_n594_n6780# a_500_n5444# 0.0023f
C70 w_n594_636# a_500_n500# 0.0023f
C71 a_500_n5444# a_n558_n5444# 0.0663f
C72 w_n594_5580# a_n500_6819# 0.00575f
C73 a_500_n7916# a_500_n6680# 0.0105f
C74 a_n558_n10388# a_n558_n9152# 0.0105f
C75 a_500_5680# w_n594_6816# 0.0023f
C76 a_n558_n7916# a_500_n7916# 0.0663f
C77 w_n594_6816# a_n500_8055# 0.00575f
C78 w_n594_n4308# a_n558_n2972# 0.0023f
C79 a_n500_639# w_n594_n600# 0.00575f
C80 a_n558_n2972# a_500_n2972# 0.0663f
C81 w_n594_n1836# a_500_n500# 0.0023f
C82 w_n594_n1836# a_n500_n3069# 0.00575f
C83 a_500_n10388# w_n594_n9252# 0.0023f
C84 a_n558_n4208# a_500_n4208# 0.0663f
C85 a_n558_3208# w_n594_1872# 0.0023f
C86 a_500_8152# w_n594_9288# 0.0023f
C87 a_n558_n7916# a_n500_n8013# 0.204f
C88 a_500_736# a_500_n500# 0.0105f
C89 w_n594_n6780# a_500_n6680# 0.0187f
C90 w_n594_n6780# a_n558_n7916# 0.0023f
C91 a_n500_n10485# w_n594_n9252# 0.00575f
C92 a_n500_5583# w_n594_4344# 0.00575f
C93 a_n558_736# a_n558_n500# 0.0105f
C94 w_n594_n8016# a_n500_n9249# 0.00575f
C95 a_n558_4444# a_n558_3208# 0.0105f
C96 w_n594_6816# a_n558_6916# 0.0187f
C97 a_500_3208# w_n594_1872# 0.0023f
C98 w_n594_1872# a_n500_1875# 0.593f
C99 a_n500_4347# w_n594_4344# 0.593f
C100 a_n500_5583# a_n500_6819# 1.03f
C101 a_500_n6680# a_n500_n6777# 0.204f
C102 a_n558_9388# a_500_9388# 0.0663f
C103 a_n558_n1736# a_n558_n500# 0.0105f
C104 a_500_6916# w_n594_5580# 0.0023f
C105 a_n500_639# a_n500_1875# 1.03f
C106 a_500_8152# a_n558_8152# 0.0663f
C107 a_n500_n4305# a_n500_n3069# 1.03f
C108 w_n594_n3072# a_n558_n1736# 0.0023f
C109 w_n594_n8016# a_500_n7916# 0.0187f
C110 w_n594_636# a_500_736# 0.0187f
C111 a_n500_n597# a_n500_639# 1.03f
C112 a_n558_n1736# a_n500_n1833# 0.204f
C113 a_n558_4444# a_n558_5680# 0.0105f
C114 a_n558_736# w_n594_n600# 0.0023f
C115 a_500_n10388# a_n558_n10388# 0.0663f
C116 a_n500_n10485# a_n500_n9249# 1.03f
C117 w_n594_n8016# a_n500_n8013# 0.593f
C118 w_n594_n4308# a_n558_n5444# 0.0023f
C119 w_n594_3108# a_n500_3111# 0.593f
C120 w_n594_8052# a_n558_8152# 0.0187f
C121 w_n594_n5544# a_n500_n4305# 0.00575f
C122 a_n558_n1736# w_n594_n600# 0.0023f
C123 w_n594_1872# a_n500_639# 0.00575f
C124 a_n558_n10388# a_n500_n10485# 0.204f
C125 w_n594_5580# a_n558_5680# 0.0187f
C126 w_n594_n10488# a_n500_n9249# 0.00575f
C127 a_500_n4208# a_500_n5444# 0.0105f
C128 w_n594_n6780# a_n500_n5541# 0.00575f
C129 a_n500_9291# a_n500_8055# 1.03f
C130 w_n594_n3072# a_500_n2972# 0.0187f
C131 a_n558_n2972# a_n500_n3069# 0.204f
C132 a_n500_n5541# a_n558_n5444# 0.204f
C133 a_n500_9291# a_500_9388# 0.204f
C134 a_n558_1972# a_n558_3208# 0.0105f
C135 w_n594_n8016# a_n500_n6777# 0.00575f
C136 a_500_3208# a_500_1972# 0.0105f
C137 a_n558_n10388# w_n594_n10488# 0.0187f
C138 a_500_n9152# w_n594_n9252# 0.0187f
C139 a_n500_1875# a_500_1972# 0.204f
C140 w_n594_n6780# a_n558_n6680# 0.0187f
C141 a_n500_n5541# a_n500_n6777# 1.03f
C142 a_n558_n6680# a_n558_n5444# 0.0105f
C143 a_n558_1972# a_n500_1875# 0.204f
C144 a_n558_736# w_n594_1872# 0.0023f
C145 w_n594_4344# a_500_4444# 0.0187f
C146 a_n500_9291# a_n558_9388# 0.204f
C147 a_n500_n6777# a_n558_n6680# 0.204f
C148 a_n500_5583# a_n558_5680# 0.204f
C149 a_n558_736# a_n500_639# 0.204f
C150 w_n594_1872# a_500_1972# 0.0187f
C151 a_n558_4444# w_n594_5580# 0.0023f
C152 a_500_n9152# a_n500_n9249# 0.204f
C153 w_n594_n1836# a_n558_n2972# 0.0023f
C154 a_n558_n4208# w_n594_n4308# 0.0187f
C155 a_500_5680# w_n594_4344# 0.0023f
C156 a_n558_1972# w_n594_1872# 0.0187f
C157 a_500_8152# a_n500_8055# 0.204f
C158 w_n594_n3072# a_500_n1736# 0.0023f
C159 a_500_n4208# a_500_n2972# 0.0105f
C160 w_n594_n4308# a_500_n4208# 0.0187f
C161 a_500_n7916# a_500_n9152# 0.0105f
C162 a_n500_n1833# a_500_n1736# 0.204f
C163 a_500_8152# a_500_9388# 0.0105f
C164 a_500_8152# w_n594_6816# 0.0023f
C165 a_n500_8055# a_n500_6819# 1.03f
C166 a_500_n500# a_n558_n500# 0.0663f
C167 w_n594_6816# a_n500_6819# 0.593f
C168 w_n594_n5544# a_n558_n5444# 0.0187f
C169 w_n594_n3072# a_n500_n3069# 0.593f
C170 a_500_n6680# a_500_n5444# 0.0105f
C171 a_500_n1736# w_n594_n600# 0.0023f
C172 a_n500_n1833# a_n500_n3069# 1.03f
C173 w_n594_8052# a_n500_8055# 0.593f
C174 w_n594_8052# a_500_9388# 0.0023f
C175 a_n558_4444# a_n500_4347# 0.204f
C176 a_n558_6916# a_n500_6819# 0.204f
C177 w_n594_n5544# a_n500_n6777# 0.00575f
C178 a_500_n500# w_n594_n600# 0.0187f
C179 w_n594_636# a_n558_n500# 0.0023f
C180 a_n500_5583# w_n594_5580# 0.593f
C181 a_n558_3208# w_n594_3108# 0.0187f
C182 w_n594_8052# a_n558_6916# 0.0023f
C183 w_n594_n9252# a_n500_n9249# 0.593f
C184 a_n558_736# a_n558_1972# 0.0105f
C185 a_500_6916# a_500_5680# 0.0105f
C186 a_n500_4347# w_n594_5580# 0.00575f
C187 a_n558_1972# a_500_1972# 0.0663f
C188 w_n594_n1836# a_n558_n500# 0.0023f
C189 w_n594_8052# a_n558_9388# 0.0023f
C190 a_500_6916# w_n594_6816# 0.0187f
C191 w_n594_n4308# a_500_n5444# 0.0023f
C192 a_n558_n10388# w_n594_n9252# 0.0023f
C193 a_n558_n7916# a_n558_n9152# 0.0105f
C194 a_500_3208# a_500_4444# 0.0105f
C195 a_500_3208# w_n594_3108# 0.0187f
C196 w_n594_n1836# a_n500_n1833# 0.593f
C197 a_500_n7916# w_n594_n9252# 0.0023f
C198 w_n594_3108# a_n500_1875# 0.00575f
C199 a_500_6916# a_n558_6916# 0.0663f
C200 a_n500_n597# a_500_n500# 0.204f
C201 w_n594_n9252# a_n500_n8013# 0.00575f
C202 w_n594_4344# a_n500_3111# 0.00575f
C203 w_n594_9288# a_n558_8152# 0.0023f
C204 a_n500_n5541# a_500_n5444# 0.204f
C205 a_500_5680# a_n558_5680# 0.0663f
C206 a_n558_n4208# w_n594_n5544# 0.0023f
C207 a_500_736# w_n594_n600# 0.0023f
C208 a_n500_4347# a_n500_5583# 1.03f
C209 w_n594_6816# a_n558_5680# 0.0023f
C210 w_n594_n8016# a_500_n6680# 0.0023f
C211 w_n594_n3072# a_n500_n4305# 0.00575f
C212 w_n594_636# a_n500_1875# 0.00575f
C213 w_n594_n8016# a_n558_n7916# 0.0187f
C214 w_n594_n5544# a_500_n4208# 0.0023f
C215 w_n594_n8016# a_n558_n9152# 0.0023f
C216 a_n500_9291# w_n594_8052# 0.00575f
C217 w_n594_636# a_n500_n597# 0.00575f
C218 a_n558_4444# a_500_4444# 0.0663f
C219 a_n500_n8013# a_n500_n9249# 1.03f
C220 a_n558_6916# a_n558_5680# 0.0105f
C221 a_n558_4444# w_n594_3108# 0.0023f
C222 w_n594_n4308# a_500_n2972# 0.0023f
C223 w_n594_n1836# a_n500_n597# 0.00575f
C224 a_500_n6680# a_n558_n6680# 0.0663f
C225 a_500_n7916# a_n500_n8013# 0.204f
C226 a_n558_n7916# a_n558_n6680# 0.0105f
C227 w_n594_636# a_n500_639# 0.593f
C228 w_n594_5580# a_500_4444# 0.0023f
C229 w_n594_n6780# a_500_n7916# 0.0023f
C230 w_n594_n3072# a_n558_n2972# 0.0187f
C231 a_n558_n4208# a_n500_n4305# 0.204f
C232 a_n558_n1736# a_500_n1736# 0.0663f
C233 w_n594_n4308# a_n500_n5541# 0.00575f
C234 a_n558_3208# a_n500_3111# 0.204f
C235 w_n594_n6780# a_n500_n8013# 0.00575f
C236 a_500_736# w_n594_1872# 0.0023f
C237 a_500_5680# w_n594_5580# 0.0187f
C238 w_n594_3108# a_500_1972# 0.0023f
C239 w_n594_n10488# a_n558_n9152# 0.0023f
C240 a_500_n4208# a_n500_n4305# 0.204f
C241 a_500_736# a_n500_639# 0.204f
C242 w_n594_n5544# a_500_n5444# 0.0187f
C243 w_n594_n6780# a_n558_n5444# 0.0023f
C244 a_500_8152# w_n594_8052# 0.0187f
C245 a_500_3208# a_n500_3111# 0.204f
C246 a_500_n10388# VSUBS 0.561f
C247 a_n558_n10388# VSUBS 0.561f
C248 a_n500_n10485# VSUBS 1.74f
C249 a_500_n9152# VSUBS 0.548f
C250 a_n558_n9152# VSUBS 0.548f
C251 a_n500_n9249# VSUBS 1.17f
C252 a_500_n7916# VSUBS 0.548f
C253 a_n558_n7916# VSUBS 0.548f
C254 a_n500_n8013# VSUBS 1.17f
C255 a_500_n6680# VSUBS 0.548f
C256 a_n558_n6680# VSUBS 0.548f
C257 a_n500_n6777# VSUBS 1.17f
C258 a_500_n5444# VSUBS 0.548f
C259 a_n558_n5444# VSUBS 0.548f
C260 a_n500_n5541# VSUBS 1.17f
C261 a_500_n4208# VSUBS 0.548f
C262 a_n558_n4208# VSUBS 0.548f
C263 a_n500_n4305# VSUBS 1.17f
C264 a_500_n2972# VSUBS 0.548f
C265 a_n558_n2972# VSUBS 0.548f
C266 a_n500_n3069# VSUBS 1.17f
C267 a_500_n1736# VSUBS 0.548f
C268 a_n558_n1736# VSUBS 0.548f
C269 a_n500_n1833# VSUBS 1.17f
C270 a_500_n500# VSUBS 0.548f
C271 a_n558_n500# VSUBS 0.548f
C272 a_n500_n597# VSUBS 1.17f
C273 a_500_736# VSUBS 0.548f
C274 a_n558_736# VSUBS 0.548f
C275 a_n500_639# VSUBS 1.17f
C276 a_500_1972# VSUBS 0.548f
C277 a_n558_1972# VSUBS 0.548f
C278 a_n500_1875# VSUBS 1.17f
C279 a_500_3208# VSUBS 0.548f
C280 a_n558_3208# VSUBS 0.548f
C281 a_n500_3111# VSUBS 1.17f
C282 a_500_4444# VSUBS 0.548f
C283 a_n558_4444# VSUBS 0.548f
C284 a_n500_4347# VSUBS 1.17f
C285 a_500_5680# VSUBS 0.548f
C286 a_n558_5680# VSUBS 0.548f
C287 a_n500_5583# VSUBS 1.17f
C288 a_500_6916# VSUBS 0.548f
C289 a_n558_6916# VSUBS 0.548f
C290 a_n500_6819# VSUBS 1.17f
C291 a_500_8152# VSUBS 0.548f
C292 a_n558_8152# VSUBS 0.548f
C293 a_n500_8055# VSUBS 1.17f
C294 a_500_9388# VSUBS 0.561f
C295 a_n558_9388# VSUBS 0.561f
C296 a_n500_9291# VSUBS 1.74f
C297 w_n594_n10488# VSUBS 4.28f
C298 w_n594_n9252# VSUBS 4.28f
C299 w_n594_n8016# VSUBS 4.28f
C300 w_n594_n6780# VSUBS 4.28f
C301 w_n594_n5544# VSUBS 4.28f
C302 w_n594_n4308# VSUBS 4.28f
C303 w_n594_n3072# VSUBS 4.28f
C304 w_n594_n1836# VSUBS 4.28f
C305 w_n594_n600# VSUBS 4.28f
C306 w_n594_636# VSUBS 4.28f
C307 w_n594_1872# VSUBS 4.28f
C308 w_n594_3108# VSUBS 4.28f
C309 w_n594_4344# VSUBS 4.28f
C310 w_n594_5580# VSUBS 4.28f
C311 w_n594_6816# VSUBS 4.28f
C312 w_n594_8052# VSUBS 4.28f
C313 w_n594_9288# VSUBS 4.28f
.ends

.subckt sky130_fd_pr__pfet_01v8_RRU5GE a_n300_n1833# w_n394_n1836# a_n358_n1736# a_300_736#
+ w_n394_636# a_n300_n597# a_300_n500# a_n300_639# w_n394_n600# a_300_n1736# a_n358_n500#
+ a_n358_736# VSUBS
X0 a_300_n500# a_n300_n597# a_n358_n500# w_n394_n600# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=3
**devattr s=58000,2116 d=58000,2116
X1 a_300_736# a_n300_639# a_n358_736# w_n394_636# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=3
**devattr s=58000,2116 d=58000,2116
X2 a_300_n1736# a_n300_n1833# a_n358_n1736# w_n394_n1836# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=3
**devattr s=58000,2116 d=58000,2116
C0 a_300_n500# w_n394_636# 0.0023f
C1 a_n300_639# w_n394_n600# 0.00346f
C2 w_n394_636# a_n358_n500# 0.0023f
C3 a_300_n1736# a_n358_n1736# 0.107f
C4 a_300_n1736# w_n394_n1836# 0.0187f
C5 a_n300_639# w_n394_636# 0.382f
C6 a_n358_736# a_n358_n500# 0.0105f
C7 a_n358_n1736# a_n358_n500# 0.0105f
C8 w_n394_n600# a_n300_n1833# 0.00346f
C9 a_300_n500# a_300_736# 0.0105f
C10 a_300_n500# a_n300_n597# 0.184f
C11 a_300_n500# w_n394_n1836# 0.0023f
C12 a_n300_n597# a_n358_n500# 0.184f
C13 w_n394_n1836# a_n358_n500# 0.0023f
C14 a_n358_736# a_n300_639# 0.184f
C15 a_n358_736# w_n394_n600# 0.0023f
C16 a_n358_n1736# w_n394_n600# 0.0023f
C17 a_n300_639# a_300_736# 0.184f
C18 a_n300_639# a_n300_n597# 0.62f
C19 w_n394_n600# a_300_736# 0.0023f
C20 a_n300_n597# w_n394_n600# 0.382f
C21 a_n358_736# w_n394_636# 0.0187f
C22 a_n358_n1736# a_n300_n1833# 0.184f
C23 a_300_n1736# a_300_n500# 0.0105f
C24 w_n394_636# a_300_736# 0.0187f
C25 a_n300_n597# w_n394_636# 0.00346f
C26 a_n300_n597# a_n300_n1833# 0.62f
C27 w_n394_n1836# a_n300_n1833# 0.382f
C28 a_300_n500# a_n358_n500# 0.107f
C29 a_n358_736# a_300_736# 0.107f
C30 a_n358_n1736# w_n394_n1836# 0.0187f
C31 a_300_n1736# w_n394_n600# 0.0023f
C32 a_n300_n597# w_n394_n1836# 0.00346f
C33 a_300_n500# w_n394_n600# 0.0187f
C34 w_n394_n600# a_n358_n500# 0.0187f
C35 a_300_n1736# a_n300_n1833# 0.184f
C36 a_300_n1736# VSUBS 0.536f
C37 a_n358_n1736# VSUBS 0.536f
C38 a_n300_n1833# VSUBS 1.08f
C39 a_300_n500# VSUBS 0.524f
C40 a_n358_n500# VSUBS 0.524f
C41 a_n300_n597# VSUBS 0.739f
C42 a_300_736# VSUBS 0.536f
C43 a_n358_736# VSUBS 0.536f
C44 a_n300_639# VSUBS 1.08f
C45 w_n394_n1836# VSUBS 2.84f
C46 w_n394_n600# VSUBS 2.84f
C47 w_n394_636# VSUBS 2.84f
.ends

.subckt sky130_fd_pr__pfet_01v8_SLZ774 w_n1594_n600# a_n1500_n597# a_1500_n500# a_n1558_n500#
+ VSUBS
X0 a_1500_n500# a_n1500_n597# a_n1558_n500# w_n1594_n600# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
C0 w_n1594_n600# a_n1500_n597# 1.65f
C1 a_n1558_n500# w_n1594_n600# 0.0187f
C2 a_n1558_n500# a_n1500_n597# 0.217f
C3 a_1500_n500# w_n1594_n600# 0.0187f
C4 a_1500_n500# a_n1500_n597# 0.217f
C5 a_1500_n500# VSUBS 0.65f
C6 a_n1558_n500# VSUBS 0.65f
C7 a_n1500_n597# VSUBS 6.74f
C8 w_n1594_n600# VSUBS 11.5f
.ends

.subckt opamp_cascode IN_P IN_M VCC VSS OUT VB_A VB_B IB
Xsky130_fd_pr__nfet_01v8_SCE452_3 VSS bias21 bias21 VSS sky130_fd_pr__nfet_01v8_SCE452
XXM9_dummy_15 VCC bias1 dummy_9 dummy_9 VSS sky130_fd_pr__pfet_01v8_ZLZ7XS
XXM5_1 VCC IN_M IN_M bias3 VCC VCC m1_44990_37960# m1_44990_37960# m1_44990_37960#
+ bias3 IN_M bias3 m1_44990_37960# bias3 IN_M m1_44990_37960# bias3 VCC IN_M IN_M
+ bias3 VCC IN_M IN_M IN_M VCC VCC VCC IN_M IN_M IN_M m1_44990_37960# m1_44990_37960#
+ m1_44990_37960# bias3 IN_M VCC bias3 m1_44990_37960# bias3 m1_44990_37960# IN_M
+ VCC bias3 m1_44990_37960# VCC bias3 VCC VCC m1_44990_37960# bias3 m1_44990_37960#
+ bias3 bias3 m1_44990_37960# bias3 VCC m1_44990_37960# IN_M VCC VSS sky130_fd_pr__pfet_01v8_7DHACV
XXM4_dummy_2 dummy_4 bias3 dummy_4 dummy_4 bias3 dummy_4 bias3 dummy_4 bias3 dummy_4
+ dummy_4 dummy_4 dummy_4 dummy_4 bias3 dummy_4 dummy_4 bias3 VSS sky130_fd_pr__nfet_01v8_MHE452
XXM9_dummy_16 VCC bias1 dummy_9 dummy_9 VSS sky130_fd_pr__pfet_01v8_ZLZ7XS
XXM100_4 IB VCC IB IB VCC VCC VCC IB VSS sky130_fd_pr__pfet_01v8_P2UXFR
XXM4_dummy_3 dummy_4 bias3 dummy_4 VSS sky130_fd_pr__nfet_01v8_SCE452
XXM9_dummy_17 VCC bias1 dummy_9 dummy_9 VSS sky130_fd_pr__pfet_01v8_ZLZ7XS
XXM5_dummy_10 dummy_5 IN_P VCC dummy_5 VSS sky130_fd_pr__pfet_01v8_MGA63L
XXM9_dummy_18 VCC bias1 dummy_9 dummy_9 VSS sky130_fd_pr__pfet_01v8_ZLZ7XS
Xsky130_fd_pr__nfet_01v8_VT3ZQW_0 dummy_4 bias3 dummy_4 VSS sky130_fd_pr__nfet_01v8_VT3ZQW
XXM9_dummy_19 VCC bias1 dummy_9 dummy_9 VSS sky130_fd_pr__pfet_01v8_ZLZ7XS
Xsky130_fd_pr__pfet_01v8_RRUZAE_0 dummy_100 IB IB VCC VCC dummy_100 dummy_100 dummy_100
+ dummy_100 VCC VCC IB dummy_100 IB dummy_100 IB VCC dummy_100 dummy_100 dummy_100
+ VSS sky130_fd_pr__pfet_01v8_RRUZAE
Xsky130_fd_pr__pfet_01v8_P2UXFR_0 IB VCC VCC IB IB VCC IB VCC VSS sky130_fd_pr__pfet_01v8_P2UXFR
XXM4_dummy_7 dummy_4 bias3 dummy_4 VSS sky130_fd_pr__nfet_01v8_SCE452
Xsky130_fd_pr__pfet_01v8_ZLZ7XS_0 VCC bias1 dummy_9 dummy_9 VSS sky130_fd_pr__pfet_01v8_ZLZ7XS
Xsky130_fd_pr__pfet_01v8_8DHNHY_0 VCC IN_P IN_P dummy_5 IN_P VCC dummy_5 VCC dummy_5
+ dummy_5 dummy_5 dummy_5 IN_P dummy_5 dummy_5 VCC dummy_5 IN_P dummy_5 dummy_5 VCC
+ dummy_5 IN_P IN_P dummy_5 VCC IN_P IN_P IN_P VCC VCC dummy_5 VCC IN_P IN_P VCC IN_P
+ dummy_5 dummy_5 dummy_5 dummy_5 IN_P VCC dummy_5 dummy_5 dummy_5 dummy_5 IN_P VCC
+ dummy_5 dummy_5 VCC dummy_5 dummy_5 VCC VCC dummy_5 dummy_5 dummy_5 dummy_5 dummy_5
+ dummy_5 dummy_5 VCC IN_P dummy_5 IN_P VCC VSS sky130_fd_pr__pfet_01v8_8DHNHY
XXM100_dummy_1 dummy_100 IB IB VCC VCC dummy_100 dummy_100 dummy_100 dummy_100 VCC
+ VCC IB dummy_100 IB dummy_100 IB VCC dummy_100 dummy_100 dummy_100 VSS sky130_fd_pr__pfet_01v8_RRUZAE
XXM1_1 m1m2 m1m2 bias1 VCC bias1 m1m2 VCC bias1 VCC VCC VCC bias1 m1m2 VCC VCC m1m2
+ VCC bias1 bias1 VCC VCC VCC bias1 m1m2 m1m2 m1m2 m1m2 bias1 VCC m1m2 VCC bias1 VCC
+ VCC VCC m1m2 m1m2 VCC bias1 VCC bias1 m1m2 bias1 VCC m1m2 VCC bias1 m1m2 VCC bias1
+ m1m2 VCC VCC VCC VCC VCC bias1 VCC VCC bias1 m1m2 m1m2 bias1 bias1 VCC VCC VCC m1m2
+ bias1 VCC bias1 VCC m1m2 VCC bias1 m1m2 VCC VCC VCC VCC VCC m1m2 VCC m1m2 bias1
+ m1m2 bias1 VCC bias1 bias1 bias1 VCC VCC VCC bias1 m1m2 VCC m1m2 VCC bias1 m1m2
+ m1m2 VCC VCC bias1 VCC m1m2 m1m2 VCC bias1 VCC m1m2 m1m2 bias1 VCC bias1 VCC VCC
+ m1m2 m1m2 VCC bias1 VCC VCC m1m2 VCC bias1 bias1 VCC VCC m1m2 VCC bias1 m1m2 VCC
+ m1m2 bias1 VCC VCC VCC m1m2 m1m2 VCC VCC VCC VCC VCC bias1 bias1 m1m2 m1m2 VCC m1m2
+ VCC VCC m1m2 VCC VCC VCC bias1 VCC m1m2 bias1 VCC VCC m1m2 m1m2 m1m2 VCC VCC m1m2
+ VCC VCC VCC m1m2 bias1 m1m2 bias1 bias1 VCC bias1 VCC VCC bias1 VCC bias1 VCC m1m2
+ VCC m1m2 m1m2 bias1 bias1 VCC bias1 bias1 VCC bias1 VCC m1m2 m1m2 VCC bias1 bias1
+ VCC VCC m1m2 m1m2 bias1 VCC bias1 VCC VCC VCC VCC bias1 m1m2 m1m2 bias1 m1m2 bias1
+ VCC VCC VCC VCC bias1 m1m2 m1m2 VCC bias1 bias1 VCC VCC bias1 VCC VCC m1m2 bias1
+ VCC VCC VCC bias1 m1m2 bias1 VCC bias1 VCC VCC bias1 VCC VCC VCC bias1 VCC bias1
+ m1m2 m1m2 VCC VCC VCC VCC bias1 VCC VCC VCC VCC VCC m1m2 bias1 bias1 VCC m1m2 VCC
+ VCC VCC bias1 bias1 VCC VCC VCC VCC m1m2 m1m2 m1m2 VCC VCC VCC VCC bias1 VCC VCC
+ m1m2 bias1 VCC VCC VCC bias1 bias1 VCC VCC m1m2 m1m2 bias1 m1m2 VCC VCC bias1 m1m2
+ VCC bias1 m1m2 m1m2 VCC VCC m1m2 VCC VCC m1m2 VCC bias1 m1m2 m1m2 bias1 m1m2 VCC
+ bias1 VCC VCC bias1 VCC bias1 VCC VCC bias1 VCC VCC VCC m1m2 VCC VCC VCC bias1 VCC
+ m1m2 VCC bias1 m1m2 VCC m1m2 m1m2 m1m2 VCC bias1 m1m2 VCC VCC VCC VCC bias1 VCC
+ bias1 m1m2 VCC m1m2 VCC m1m2 VCC VCC VCC bias1 VCC bias1 bias1 m1m2 bias1 VCC VCC
+ VCC VCC VCC VCC VCC VCC bias1 VCC VCC m1m2 bias1 VCC VCC bias1 VCC m1m2 m1m2 VCC
+ m1m2 VCC VCC VSS VCC m1m2 sky130_fd_pr__pfet_01v8_F76D73
XXM4_dummy_9 dummy_4 bias3 dummy_4 VSS sky130_fd_pr__nfet_01v8_SCE452
XXM1_2 m1m2 m1m2 bias1 VCC bias1 m1m2 VCC bias1 VCC VCC VCC bias1 m1m2 VCC VCC m1m2
+ VCC bias1 bias1 VCC VCC VCC bias1 m1m2 m1m2 m1m2 m1m2 bias1 VCC m1m2 VCC bias1 VCC
+ VCC VCC m1m2 m1m2 VCC bias1 VCC bias1 m1m2 bias1 VCC m1m2 VCC bias1 m1m2 VCC bias1
+ m1m2 VCC VCC VCC VCC VCC bias1 VCC VCC bias1 m1m2 m1m2 bias1 bias1 VCC VCC VCC m1m2
+ bias1 VCC bias1 VCC m1m2 VCC bias1 m1m2 VCC VCC VCC VCC VCC m1m2 VCC m1m2 bias1
+ m1m2 bias1 VCC bias1 bias1 bias1 VCC VCC VCC bias1 m1m2 VCC m1m2 VCC bias1 m1m2
+ m1m2 VCC VCC bias1 VCC m1m2 m1m2 VCC bias1 VCC m1m2 m1m2 bias1 VCC bias1 VCC VCC
+ m1m2 m1m2 VCC bias1 VCC VCC m1m2 VCC bias1 bias1 VCC VCC m1m2 VCC bias1 m1m2 VCC
+ m1m2 bias1 VCC VCC VCC m1m2 m1m2 VCC VCC VCC VCC VCC bias1 bias1 m1m2 m1m2 VCC m1m2
+ VCC VCC m1m2 VCC VCC VCC bias1 VCC m1m2 bias1 VCC VCC m1m2 m1m2 m1m2 VCC VCC m1m2
+ VCC VCC VCC m1m2 bias1 m1m2 bias1 bias1 VCC bias1 VCC VCC bias1 VCC bias1 VCC m1m2
+ VCC m1m2 m1m2 bias1 bias1 VCC bias1 bias1 VCC bias1 VCC m1m2 m1m2 VCC bias1 bias1
+ VCC VCC m1m2 m1m2 bias1 VCC bias1 VCC VCC VCC VCC bias1 m1m2 m1m2 bias1 m1m2 bias1
+ VCC VCC VCC VCC bias1 m1m2 m1m2 VCC bias1 bias1 VCC VCC bias1 VCC VCC m1m2 bias1
+ VCC VCC VCC bias1 m1m2 bias1 VCC bias1 VCC VCC bias1 VCC VCC VCC bias1 VCC bias1
+ m1m2 m1m2 VCC VCC VCC VCC bias1 VCC VCC VCC VCC VCC m1m2 bias1 bias1 VCC m1m2 VCC
+ VCC VCC bias1 bias1 VCC VCC VCC VCC m1m2 m1m2 m1m2 VCC VCC VCC VCC bias1 VCC VCC
+ m1m2 bias1 VCC VCC VCC bias1 bias1 VCC VCC m1m2 m1m2 bias1 m1m2 VCC VCC bias1 m1m2
+ VCC bias1 m1m2 m1m2 VCC VCC m1m2 VCC VCC m1m2 VCC bias1 m1m2 m1m2 bias1 m1m2 VCC
+ bias1 VCC VCC bias1 VCC bias1 VCC VCC bias1 VCC VCC VCC m1m2 VCC VCC VCC bias1 VCC
+ m1m2 VCC bias1 m1m2 VCC m1m2 m1m2 m1m2 VCC bias1 m1m2 VCC VCC VCC VCC bias1 VCC
+ bias1 m1m2 VCC m1m2 VCC m1m2 VCC VCC VCC bias1 VCC bias1 bias1 m1m2 bias1 VCC VCC
+ VCC VCC VCC VCC VCC VCC bias1 VCC VCC m1m2 bias1 VCC VCC bias1 VCC m1m2 m1m2 VCC
+ m1m2 VCC VCC VSS VCC m1m2 sky130_fd_pr__pfet_01v8_F76D73
XXM3_dummy_1 VB_B dummy_3 dummy_3 dummy_3 VB_B dummy_3 VB_B VB_B VB_B VB_B dummy_3
+ dummy_3 dummy_3 dummy_3 dummy_3 dummy_3 VB_B dummy_3 dummy_3 dummy_3 VB_B dummy_3
+ dummy_3 dummy_3 VB_B dummy_3 dummy_3 dummy_3 dummy_3 VB_B dummy_3 dummy_3 VB_B VB_B
+ dummy_3 dummy_3 VB_B dummy_3 VB_B dummy_3 VB_B VB_B dummy_3 VB_B dummy_3 dummy_3
+ dummy_3 dummy_3 dummy_3 dummy_3 dummy_3 VSS sky130_fd_pr__nfet_01v8_WK8VRD
XXM100_dummy_3 IB VCC dummy_100 IB dummy_100 VCC dummy_100 dummy_100 VSS sky130_fd_pr__pfet_01v8_P2UXFR
XXM1_3 m1m2 m1m2 bias1 VCC bias1 m1m2 VCC bias1 VCC VCC VCC bias1 m1m2 VCC VCC m1m2
+ VCC bias1 bias1 VCC VCC VCC bias1 m1m2 m1m2 m1m2 m1m2 bias1 VCC m1m2 VCC bias1 VCC
+ VCC VCC m1m2 m1m2 VCC bias1 VCC bias1 m1m2 bias1 VCC m1m2 VCC bias1 m1m2 VCC bias1
+ m1m2 VCC VCC VCC VCC VCC bias1 VCC VCC bias1 m1m2 m1m2 bias1 bias1 VCC VCC VCC m1m2
+ bias1 VCC bias1 VCC m1m2 VCC bias1 m1m2 VCC VCC VCC VCC VCC m1m2 VCC m1m2 bias1
+ m1m2 bias1 VCC bias1 bias1 bias1 VCC VCC VCC bias1 m1m2 VCC m1m2 VCC bias1 m1m2
+ m1m2 VCC VCC bias1 VCC m1m2 m1m2 VCC bias1 VCC m1m2 m1m2 bias1 VCC bias1 VCC VCC
+ m1m2 m1m2 VCC bias1 VCC VCC m1m2 VCC bias1 bias1 VCC VCC m1m2 VCC bias1 m1m2 VCC
+ m1m2 bias1 VCC VCC VCC m1m2 m1m2 VCC VCC VCC VCC VCC bias1 bias1 m1m2 m1m2 VCC m1m2
+ VCC VCC m1m2 VCC VCC VCC bias1 VCC m1m2 bias1 VCC VCC m1m2 m1m2 m1m2 VCC VCC m1m2
+ VCC VCC VCC m1m2 bias1 m1m2 bias1 bias1 VCC bias1 VCC VCC bias1 VCC bias1 VCC m1m2
+ VCC m1m2 m1m2 bias1 bias1 VCC bias1 bias1 VCC bias1 VCC m1m2 m1m2 VCC bias1 bias1
+ VCC VCC m1m2 m1m2 bias1 VCC bias1 VCC VCC VCC VCC bias1 m1m2 m1m2 bias1 m1m2 bias1
+ VCC VCC VCC VCC bias1 m1m2 m1m2 VCC bias1 bias1 VCC VCC bias1 VCC VCC m1m2 bias1
+ VCC VCC VCC bias1 m1m2 bias1 VCC bias1 VCC VCC bias1 VCC VCC VCC bias1 VCC bias1
+ m1m2 m1m2 VCC VCC VCC VCC bias1 VCC VCC VCC VCC VCC m1m2 bias1 bias1 VCC m1m2 VCC
+ VCC VCC bias1 bias1 VCC VCC VCC VCC m1m2 m1m2 m1m2 VCC VCC VCC VCC bias1 VCC VCC
+ m1m2 bias1 VCC VCC VCC bias1 bias1 VCC VCC m1m2 m1m2 bias1 m1m2 VCC VCC bias1 m1m2
+ VCC bias1 m1m2 m1m2 VCC VCC m1m2 VCC VCC m1m2 VCC bias1 m1m2 m1m2 bias1 m1m2 VCC
+ bias1 VCC VCC bias1 VCC bias1 VCC VCC bias1 VCC VCC VCC m1m2 VCC VCC VCC bias1 VCC
+ m1m2 VCC bias1 m1m2 VCC m1m2 m1m2 m1m2 VCC bias1 m1m2 VCC VCC VCC VCC bias1 VCC
+ bias1 m1m2 VCC m1m2 VCC m1m2 VCC VCC VCC bias1 VCC bias1 bias1 m1m2 bias1 VCC VCC
+ VCC VCC VCC VCC VCC VCC bias1 VCC VCC m1m2 bias1 VCC VCC bias1 VCC m1m2 m1m2 VCC
+ m1m2 VCC VCC VSS VCC m1m2 sky130_fd_pr__pfet_01v8_F76D73
XXM100_dummy_4 IB VCC dummy_100 IB dummy_100 VCC dummy_100 dummy_100 VSS sky130_fd_pr__pfet_01v8_P2UXFR
Xsky130_fd_pr__pfet_01v8_MGA63L_0 dummy_5 IN_P VCC dummy_5 VSS sky130_fd_pr__pfet_01v8_MGA63L
XXM3_dummy_3 dummy_3 dummy_3 VB_B VSS sky130_fd_pr__nfet_01v8_AH5E2K
XXM100_dummy_5 IB dummy_100 VCC dummy_100 VSS sky130_fd_pr__pfet_01v8_C2U9V5
XXM1 m1m2 m1m2 bias1 VCC bias1 m1m2 VCC bias1 VCC VCC VCC bias1 m1m2 VCC VCC m1m2
+ VCC bias1 bias1 VCC VCC VCC bias1 m1m2 m1m2 m1m2 m1m2 bias1 VCC m1m2 VCC bias1 VCC
+ VCC VCC m1m2 m1m2 VCC bias1 VCC bias1 m1m2 bias1 VCC m1m2 VCC bias1 m1m2 VCC bias1
+ m1m2 VCC VCC VCC VCC VCC bias1 VCC VCC bias1 m1m2 m1m2 bias1 bias1 VCC VCC VCC m1m2
+ bias1 VCC bias1 VCC m1m2 VCC bias1 m1m2 VCC VCC VCC VCC VCC m1m2 VCC m1m2 bias1
+ m1m2 bias1 VCC bias1 bias1 bias1 VCC VCC VCC bias1 m1m2 VCC m1m2 VCC bias1 m1m2
+ m1m2 VCC VCC bias1 VCC m1m2 m1m2 VCC bias1 VCC m1m2 m1m2 bias1 VCC bias1 VCC VCC
+ m1m2 m1m2 VCC bias1 VCC VCC m1m2 VCC bias1 bias1 VCC VCC m1m2 VCC bias1 m1m2 VCC
+ m1m2 bias1 VCC VCC VCC m1m2 m1m2 VCC VCC VCC VCC VCC bias1 bias1 m1m2 m1m2 VCC m1m2
+ VCC VCC m1m2 VCC VCC VCC bias1 VCC m1m2 bias1 VCC VCC m1m2 m1m2 m1m2 VCC VCC m1m2
+ VCC VCC VCC m1m2 bias1 m1m2 bias1 bias1 VCC bias1 VCC VCC bias1 VCC bias1 VCC m1m2
+ VCC m1m2 m1m2 bias1 bias1 VCC bias1 bias1 VCC bias1 VCC m1m2 m1m2 VCC bias1 bias1
+ VCC VCC m1m2 m1m2 bias1 VCC bias1 VCC VCC VCC VCC bias1 m1m2 m1m2 bias1 m1m2 bias1
+ VCC VCC VCC VCC bias1 m1m2 m1m2 VCC bias1 bias1 VCC VCC bias1 VCC VCC m1m2 bias1
+ VCC VCC VCC bias1 m1m2 bias1 VCC bias1 VCC VCC bias1 VCC VCC VCC bias1 VCC bias1
+ m1m2 m1m2 VCC VCC VCC VCC bias1 VCC VCC VCC VCC VCC m1m2 bias1 bias1 VCC m1m2 VCC
+ VCC VCC bias1 bias1 VCC VCC VCC VCC m1m2 m1m2 m1m2 VCC VCC VCC VCC bias1 VCC VCC
+ m1m2 bias1 VCC VCC VCC bias1 bias1 VCC VCC m1m2 m1m2 bias1 m1m2 VCC VCC bias1 m1m2
+ VCC bias1 m1m2 m1m2 VCC VCC m1m2 VCC VCC m1m2 VCC bias1 m1m2 m1m2 bias1 m1m2 VCC
+ bias1 VCC VCC bias1 VCC bias1 VCC VCC bias1 VCC VCC VCC m1m2 VCC VCC VCC bias1 VCC
+ m1m2 VCC bias1 m1m2 VCC m1m2 m1m2 m1m2 VCC bias1 m1m2 VCC VCC VCC VCC bias1 VCC
+ bias1 m1m2 VCC m1m2 VCC m1m2 VCC VCC VCC bias1 VCC bias1 bias1 m1m2 bias1 VCC VCC
+ VCC VCC VCC VCC VCC VCC bias1 VCC VCC m1m2 bias1 VCC VCC bias1 VCC m1m2 m1m2 VCC
+ m1m2 VCC VCC VSS VCC m1m2 sky130_fd_pr__pfet_01v8_F76D73
XXM100_dummy_6 IB dummy_100 VCC dummy_100 VSS sky130_fd_pr__pfet_01v8_C2U9V5
XXM3_dummy_4 dummy_3 dummy_3 VB_B VSS sky130_fd_pr__nfet_01v8_AH5E2K
Xsky130_fd_pr__nfet_01v8_QP5WRD_0 bias1 bias1 VB_B bias1 VB_B VB_B VB_B VB_B m3m4
+ m3m4 m3m4 m3m4 bias1 bias1 VB_B bias1 bias1 VB_B bias1 bias1 m3m4 VB_B m3m4 m3m4
+ m3m4 m3m4 m3m4 VB_B VB_B bias1 bias1 VB_B bias1 VB_B bias1 VB_B VB_B m3m4 VB_B m3m4
+ m3m4 m3m4 m3m4 bias1 bias1 VSS sky130_fd_pr__nfet_01v8_QP5WRD
XXM2 bias1 VB_A m1m2 bias1 VB_A m1m2 VCC VCC m1m2 m1m2 m1m2 VB_A VCC m1m2 VCC bias1
+ VCC VCC VB_A bias1 VCC VB_A bias1 bias1 VB_A VB_A m1m2 VB_A m1m2 m1m2 bias1 m1m2
+ VCC m1m2 VCC VCC bias1 bias1 VCC bias1 bias1 bias1 VB_A VB_A VB_A VCC m1m2 VB_A
+ VCC VB_A m1m2 VCC VB_A m1m2 VCC VB_A m1m2 bias1 bias1 bias1 VSS sky130_fd_pr__pfet_01v8_UDM5A5
XXM100_dummy_7 IB dummy_100 VCC dummy_100 VSS sky130_fd_pr__pfet_01v8_C2U9V5
XXM4_dummy_10 dummy_4 bias3 dummy_4 VSS sky130_fd_pr__nfet_01v8_SCE452
XXM3 m3m4 m3m4 VB_B m3m4 VB_B VB_B VB_B VB_B bias1 bias1 bias1 bias1 m3m4 m3m4 VB_B
+ m3m4 m3m4 VB_B m3m4 m3m4 bias1 VB_B bias1 bias1 bias1 bias1 bias1 VB_B VB_B m3m4
+ m3m4 VB_B m3m4 VB_B m3m4 VB_B VB_B bias1 VB_B bias1 bias1 bias1 bias1 m3m4 m3m4
+ VSS sky130_fd_pr__nfet_01v8_QP5WRD
XXM8_1 VSS bias21 bias21 VSS sky130_fd_pr__nfet_01v8_VT3ZQW
XXM3_dummy_6 dummy_3 dummy_3 VB_B VSS sky130_fd_pr__nfet_01v8_AH5E2K
XXM100_dummy_8 IB dummy_100 VCC dummy_100 VSS sky130_fd_pr__pfet_01v8_C2U9V5
XXM4 VSS m3m4 bias3 VSS sky130_fd_pr__nfet_01v8_3ZAA45
XXM100_dummy_9 IB dummy_100 VCC dummy_100 VSS sky130_fd_pr__pfet_01v8_C2U9V5
XXM3_dummy_7 dummy_3 dummy_3 VB_B VSS sky130_fd_pr__nfet_01v8_AH5E2K
XXM5 VCC IN_M IN_M m1_44990_37960# VCC VCC bias3 bias3 bias3 m1_44990_37960# IN_M
+ m1_44990_37960# bias3 m1_44990_37960# IN_M bias3 m1_44990_37960# VCC IN_M IN_M m1_44990_37960#
+ VCC IN_M IN_M IN_M VCC VCC VCC IN_M IN_M IN_M bias3 bias3 bias3 m1_44990_37960#
+ IN_M VCC m1_44990_37960# bias3 m1_44990_37960# bias3 IN_M VCC m1_44990_37960# bias3
+ VCC m1_44990_37960# VCC VCC bias3 m1_44990_37960# bias3 m1_44990_37960# m1_44990_37960#
+ bias3 m1_44990_37960# VCC bias3 IN_M VCC VSS sky130_fd_pr__pfet_01v8_7DHACV
XXM8_3 VSS bias21 bias21 VSS sky130_fd_pr__nfet_01v8_VT3ZQW
XXM3_dummy_8 dummy_3 dummy_3 VB_B VSS sky130_fd_pr__nfet_01v8_AH5E2K
XXM6 bias3 bias3 VSS VSS sky130_fd_pr__nfet_01v8_VT3ZQW
XXM3_dummy_9 dummy_3 dummy_3 VB_B VSS sky130_fd_pr__nfet_01v8_AH5E2K
Xsky130_fd_pr__pfet_01v8_SKU9VM_0 VB_A dummy_2 VCC dummy_2 VSS sky130_fd_pr__pfet_01v8_SKU9VM
XXM6_1 bias3 bias3 VSS VSS sky130_fd_pr__nfet_01v8_VT3ZQW
XXM7 VCC IN_P IN_P bias21 VCC VCC m1_44990_37960# m1_44990_37960# m1_44990_37960#
+ bias21 IN_P bias21 m1_44990_37960# bias21 IN_P m1_44990_37960# bias21 VCC IN_P IN_P
+ bias21 VCC IN_P IN_P IN_P VCC VCC VCC IN_P IN_P IN_P m1_44990_37960# m1_44990_37960#
+ m1_44990_37960# bias21 IN_P VCC bias21 m1_44990_37960# bias21 m1_44990_37960# IN_P
+ VCC bias21 m1_44990_37960# VCC bias21 VCC VCC m1_44990_37960# bias21 m1_44990_37960#
+ bias21 bias21 m1_44990_37960# bias21 VCC m1_44990_37960# IN_P VCC VSS sky130_fd_pr__pfet_01v8_7DHACV
Xsky130_fd_pr__pfet_01v8_E769TZ_0 dummy_9 dummy_9 bias1 VCC bias1 dummy_9 dummy_9
+ bias1 VCC VCC dummy_9 bias1 dummy_9 VCC VCC dummy_9 dummy_9 dummy_9 bias1 bias1
+ VCC VCC dummy_9 bias1 dummy_9 dummy_9 dummy_9 dummy_9 bias1 VCC dummy_9 dummy_9
+ bias1 VCC dummy_9 dummy_9 dummy_9 dummy_9 VCC bias1 VCC bias1 dummy_9 bias1 dummy_9
+ dummy_9 dummy_9 bias1 dummy_9 dummy_9 bias1 dummy_9 bias1 VCC VCC dummy_9 VCC VCC
+ bias1 dummy_9 dummy_9 bias1 dummy_9 dummy_9 bias1 bias1 VCC VCC dummy_9 dummy_9
+ bias1 dummy_9 bias1 dummy_9 dummy_9 dummy_9 bias1 dummy_9 VCC VCC dummy_9 VCC VCC
+ dummy_9 VCC dummy_9 bias1 dummy_9 bias1 dummy_9 bias1 bias1 bias1 VCC dummy_9 VCC
+ bias1 dummy_9 dummy_9 dummy_9 dummy_9 bias1 dummy_9 dummy_9 VCC bias1 VCC VCC dummy_9
+ dummy_9 dummy_9 bias1 dummy_9 dummy_9 dummy_9 bias1 VCC bias1 dummy_9 VCC dummy_9
+ dummy_9 dummy_9 VCC bias1 VCC dummy_9 dummy_9 dummy_9 bias1 bias1 dummy_9 dummy_9
+ dummy_9 dummy_9 VCC bias1 dummy_9 VCC dummy_9 bias1 VCC dummy_9 VCC dummy_9 dummy_9
+ dummy_9 VCC VCC dummy_9 VCC VCC bias1 bias1 dummy_9 dummy_9 dummy_9 dummy_9 dummy_9
+ dummy_9 dummy_9 VCC VCC dummy_9 dummy_9 bias1 dummy_9 dummy_9 bias1 VCC dummy_9
+ dummy_9 dummy_9 dummy_9 VCC dummy_9 dummy_9 dummy_9 VCC VCC dummy_9 bias1 dummy_9
+ bias1 bias1 dummy_9 bias1 VCC dummy_9 bias1 VCC bias1 VCC dummy_9 VCC dummy_9 dummy_9
+ bias1 bias1 dummy_9 bias1 bias1 VCC bias1 dummy_9 dummy_9 dummy_9 VCC bias1 bias1
+ VCC VCC dummy_9 dummy_9 bias1 dummy_9 bias1 dummy_9 dummy_9 VCC bias1 dummy_9 bias1
+ dummy_9 dummy_9 bias1 dummy_9 bias1 VCC dummy_9 dummy_9 dummy_9 bias1 dummy_9 dummy_9
+ dummy_9 bias1 bias1 dummy_9 dummy_9 bias1 VCC dummy_9 dummy_9 bias1 VCC VCC dummy_9
+ bias1 dummy_9 bias1 dummy_9 bias1 VCC dummy_9 bias1 VCC dummy_9 dummy_9 bias1 dummy_9
+ bias1 dummy_9 dummy_9 VCC VCC VCC dummy_9 bias1 VCC VCC VCC dummy_9 dummy_9 dummy_9
+ bias1 bias1 dummy_9 dummy_9 VCC VCC VCC bias1 bias1 dummy_9 dummy_9 VCC VCC dummy_9
+ dummy_9 dummy_9 VCC VCC VCC VCC bias1 VCC VCC dummy_9 bias1 dummy_9 dummy_9 dummy_9
+ bias1 bias1 dummy_9 dummy_9 dummy_9 dummy_9 bias1 dummy_9 VCC VCC dummy_9 bias1
+ dummy_9 dummy_9 bias1 dummy_9 dummy_9 VCC VCC dummy_9 dummy_9 VCC dummy_9 dummy_9
+ bias1 dummy_9 dummy_9 bias1 dummy_9 dummy_9 bias1 dummy_9 VCC bias1 dummy_9 bias1
+ VCC dummy_9 bias1 VCC dummy_9 dummy_9 dummy_9 VCC VCC dummy_9 bias1 VCC dummy_9
+ dummy_9 bias1 dummy_9 VCC dummy_9 dummy_9 dummy_9 VCC bias1 dummy_9 dummy_9 VCC
+ VCC dummy_9 bias1 dummy_9 bias1 dummy_9 dummy_9 dummy_9 dummy_9 dummy_9 VCC VCC
+ dummy_9 bias1 dummy_9 bias1 bias1 dummy_9 bias1 dummy_9 dummy_9 VCC VCC VCC dummy_9
+ dummy_9 dummy_9 bias1 dummy_9 dummy_9 dummy_9 bias1 VCC VCC bias1 dummy_9 dummy_9
+ dummy_9 VCC dummy_9 VCC VCC VSS dummy_9 dummy_9 sky130_fd_pr__pfet_01v8_E769TZ
XXM6_2 bias3 bias3 VSS VSS sky130_fd_pr__nfet_01v8_VT3ZQW
XXM8 VSS bias21 bias21 VSS sky130_fd_pr__nfet_01v8_VT3ZQW
XXM2_dummy_2 dummy_2 dummy_2 VB_A VB_A dummy_2 dummy_2 VB_A dummy_2 VCC VCC dummy_2
+ dummy_2 dummy_2 VB_A VCC dummy_2 dummy_2 VCC dummy_2 VCC VCC VB_A dummy_2 VCC VB_A
+ dummy_2 VCC dummy_2 VB_A VB_A dummy_2 VB_A dummy_2 dummy_2 dummy_2 dummy_2 dummy_2
+ VCC dummy_2 VCC VCC dummy_2 dummy_2 VCC dummy_2 dummy_2 dummy_2 VB_A VB_A VB_A VCC
+ dummy_2 VB_A VB_A VCC VB_A dummy_2 VCC VB_A dummy_2 VCC dummy_2 VB_A dummy_2 dummy_2
+ VCC dummy_2 dummy_2 VSS sky130_fd_pr__pfet_01v8_UDMRD5
Xsky130_fd_pr__pfet_01v8_RRU5GE_0 IB VCC m1_44990_37960# VCC VCC IB VCC IB VCC VCC
+ m1_44990_37960# m1_44990_37960# VSS sky130_fd_pr__pfet_01v8_RRU5GE
XXM6_3 bias3 bias3 VSS VSS sky130_fd_pr__nfet_01v8_VT3ZQW
XXM9 VCC VCC bias1 VCC bias1 VCC m9m10 bias1 VCC VCC m9m10 bias1 VCC VCC m9m10 VCC
+ m9m10 bias1 bias1 VCC VCC m9m10 bias1 VCC VCC VCC VCC bias1 VCC VCC m9m10 bias1
+ VCC m9m10 m9m10 VCC VCC VCC bias1 VCC bias1 VCC bias1 m9m10 VCC m9m10 bias1 VCC
+ m9m10 bias1 VCC VCC VCC m9m10 VCC VCC bias1 m9m10 m9m10 bias1 VCC VCC bias1 bias1
+ VCC VCC m9m10 VCC bias1 m9m10 bias1 m9m10 VCC m9m10 bias1 VCC VCC VCC m9m10 VCC
+ VCC VCC VCC VCC bias1 VCC bias1 m9m10 bias1 bias1 bias1 VCC m9m10 VCC bias1 VCC
+ m9m10 VCC m9m10 bias1 VCC VCC VCC VCC bias1 VCC VCC VCC m9m10 bias1 m9m10 VCC VCC
+ bias1 VCC bias1 m9m10 VCC VCC VCC VCC bias1 VCC m9m10 VCC m9m10 bias1 bias1 m9m10
+ m9m10 VCC VCC bias1 VCC VCC VCC bias1 VCC m9m10 m9m10 VCC VCC VCC VCC m9m10 VCC
+ VCC bias1 bias1 VCC VCC m9m10 VCC m9m10 m9m10 VCC VCC VCC m9m10 bias1 m9m10 VCC
+ bias1 VCC m9m10 VCC VCC VCC VCC m9m10 VCC m9m10 VCC VCC VCC bias1 VCC bias1 bias1
+ m9m10 bias1 VCC m9m10 bias1 VCC bias1 VCC VCC VCC VCC VCC bias1 bias1 m9m10 bias1
+ bias1 VCC bias1 m9m10 VCC VCC VCC bias1 bias1 VCC VCC VCC VCC bias1 m9m10 bias1
+ m9m10 m9m10 VCC m9m10 bias1 VCC VCC bias1 VCC bias1 VCC m9m10 m9m10 m9m10 bias1
+ VCC VCC m9m10 bias1 bias1 m9m10 m9m10 bias1 VCC m9m10 VCC bias1 VCC VCC m9m10 bias1
+ VCC bias1 m9m10 bias1 VCC m9m10 bias1 VCC m9m10 m9m10 bias1 m9m10 bias1 VCC VCC
+ VCC VCC VCC m9m10 bias1 VCC VCC VCC m9m10 m9m10 VCC bias1 bias1 m9m10 VCC VCC VCC
+ VCC bias1 bias1 m9m10 m9m10 VCC VCC VCC VCC VCC VCC VCC VCC VCC bias1 VCC VCC VCC
+ bias1 m9m10 m9m10 m9m10 bias1 bias1 m9m10 m9m10 VCC VCC bias1 VCC VCC VCC bias1
+ VCC m9m10 bias1 VCC VCC VCC VCC VCC m9m10 VCC VCC m9m10 bias1 VCC VCC bias1 VCC
+ m9m10 bias1 m9m10 VCC bias1 m9m10 bias1 VCC m9m10 bias1 VCC m9m10 m9m10 VCC VCC
+ VCC m9m10 bias1 VCC VCC m9m10 bias1 VCC VCC VCC VCC VCC VCC bias1 VCC m9m10 VCC
+ VCC m9m10 bias1 m9m10 bias1 VCC m9m10 VCC m9m10 VCC VCC VCC m9m10 bias1 m9m10 bias1
+ bias1 VCC bias1 m9m10 m9m10 VCC VCC VCC m9m10 m9m10 m9m10 bias1 m9m10 m9m10 VCC
+ bias1 VCC VCC bias1 m9m10 VCC VCC VCC VCC VCC VCC VSS m9m10 VCC sky130_fd_pr__pfet_01v8_F76D73
XXM2_dummy_3 VB_A dummy_2 VCC dummy_2 VSS sky130_fd_pr__pfet_01v8_SKU9VM
Xsky130_fd_pr__pfet_01v8_C2U9V5_0 IB dummy_100 VCC dummy_100 VSS sky130_fd_pr__pfet_01v8_C2U9V5
XXM2_dummy_4 VB_A dummy_2 VCC dummy_2 VSS sky130_fd_pr__pfet_01v8_SKU9VM
XXM2_dummy_5 VB_A dummy_2 VCC dummy_2 VSS sky130_fd_pr__pfet_01v8_SKU9VM
Xsky130_fd_pr__nfet_01v8_AH5E2K_0 dummy_3 dummy_3 VB_B VSS sky130_fd_pr__nfet_01v8_AH5E2K
XXM2_1 m1m2 VB_A bias1 m1m2 VB_A bias1 VCC VCC bias1 bias1 bias1 VB_A VCC bias1 VCC
+ m1m2 VCC VCC VB_A m1m2 VCC VB_A m1m2 m1m2 VB_A VB_A bias1 VB_A bias1 bias1 m1m2
+ bias1 VCC bias1 VCC VCC m1m2 m1m2 VCC m1m2 m1m2 m1m2 VB_A VB_A VB_A VCC bias1 VB_A
+ VCC VB_A bias1 VCC VB_A bias1 VCC VB_A bias1 m1m2 m1m2 m1m2 VSS sky130_fd_pr__pfet_01v8_UDM5A5
XXM2_dummy_6 VB_A dummy_2 VCC dummy_2 VSS sky130_fd_pr__pfet_01v8_SKU9VM
Xsky130_fd_pr__nfet_01v8_3ZAA45_0 m11m12 VSS bias21 VSS sky130_fd_pr__nfet_01v8_3ZAA45
XXM3_dummy_10 dummy_3 dummy_3 VB_B VSS sky130_fd_pr__nfet_01v8_AH5E2K
Xsky130_fd_pr__nfet_01v8_MHE452_0 dummy_4 bias3 dummy_4 dummy_4 bias3 dummy_4 bias3
+ dummy_4 bias3 dummy_4 dummy_4 dummy_4 dummy_4 dummy_4 bias3 dummy_4 dummy_4 bias3
+ VSS sky130_fd_pr__nfet_01v8_MHE452
XXM2_dummy_7 VB_A dummy_2 VCC dummy_2 VSS sky130_fd_pr__pfet_01v8_SKU9VM
Xsky130_fd_pr__pfet_01v8_F76D73_0 m1m2 m1m2 bias1 VCC bias1 m1m2 VCC bias1 VCC VCC
+ VCC bias1 m1m2 VCC VCC m1m2 VCC bias1 bias1 VCC VCC VCC bias1 m1m2 m1m2 m1m2 m1m2
+ bias1 VCC m1m2 VCC bias1 VCC VCC VCC m1m2 m1m2 VCC bias1 VCC bias1 m1m2 bias1 VCC
+ m1m2 VCC bias1 m1m2 VCC bias1 m1m2 VCC VCC VCC VCC VCC bias1 VCC VCC bias1 m1m2
+ m1m2 bias1 bias1 VCC VCC VCC m1m2 bias1 VCC bias1 VCC m1m2 VCC bias1 m1m2 VCC VCC
+ VCC VCC VCC m1m2 VCC m1m2 bias1 m1m2 bias1 VCC bias1 bias1 bias1 VCC VCC VCC bias1
+ m1m2 VCC m1m2 VCC bias1 m1m2 m1m2 VCC VCC bias1 VCC m1m2 m1m2 VCC bias1 VCC m1m2
+ m1m2 bias1 VCC bias1 VCC VCC m1m2 m1m2 VCC bias1 VCC VCC m1m2 VCC bias1 bias1 VCC
+ VCC m1m2 VCC bias1 m1m2 VCC m1m2 bias1 VCC VCC VCC m1m2 m1m2 VCC VCC VCC VCC VCC
+ bias1 bias1 m1m2 m1m2 VCC m1m2 VCC VCC m1m2 VCC VCC VCC bias1 VCC m1m2 bias1 VCC
+ VCC m1m2 m1m2 m1m2 VCC VCC m1m2 VCC VCC VCC m1m2 bias1 m1m2 bias1 bias1 VCC bias1
+ VCC VCC bias1 VCC bias1 VCC m1m2 VCC m1m2 m1m2 bias1 bias1 VCC bias1 bias1 VCC bias1
+ VCC m1m2 m1m2 VCC bias1 bias1 VCC VCC m1m2 m1m2 bias1 VCC bias1 VCC VCC VCC VCC
+ bias1 m1m2 m1m2 bias1 m1m2 bias1 VCC VCC VCC VCC bias1 m1m2 m1m2 VCC bias1 bias1
+ VCC VCC bias1 VCC VCC m1m2 bias1 VCC VCC VCC bias1 m1m2 bias1 VCC bias1 VCC VCC
+ bias1 VCC VCC VCC bias1 VCC bias1 m1m2 m1m2 VCC VCC VCC VCC bias1 VCC VCC VCC VCC
+ VCC m1m2 bias1 bias1 VCC m1m2 VCC VCC VCC bias1 bias1 VCC VCC VCC VCC m1m2 m1m2
+ m1m2 VCC VCC VCC VCC bias1 VCC VCC m1m2 bias1 VCC VCC VCC bias1 bias1 VCC VCC m1m2
+ m1m2 bias1 m1m2 VCC VCC bias1 m1m2 VCC bias1 m1m2 m1m2 VCC VCC m1m2 VCC VCC m1m2
+ VCC bias1 m1m2 m1m2 bias1 m1m2 VCC bias1 VCC VCC bias1 VCC bias1 VCC VCC bias1 VCC
+ VCC VCC m1m2 VCC VCC VCC bias1 VCC m1m2 VCC bias1 m1m2 VCC m1m2 m1m2 m1m2 VCC bias1
+ m1m2 VCC VCC VCC VCC bias1 VCC bias1 m1m2 VCC m1m2 VCC m1m2 VCC VCC VCC bias1 VCC
+ bias1 bias1 m1m2 bias1 VCC VCC VCC VCC VCC VCC VCC VCC bias1 VCC VCC m1m2 bias1
+ VCC VCC bias1 VCC m1m2 m1m2 VCC m1m2 VCC VCC VSS VCC m1m2 sky130_fd_pr__pfet_01v8_F76D73
Xsky130_fd_pr__pfet_01v8_UDM5A5_0 m9m10 VB_A OUT m9m10 VB_A OUT VCC VCC OUT OUT OUT
+ VB_A VCC OUT VCC m9m10 VCC VCC VB_A m9m10 VCC VB_A m9m10 m9m10 VB_A VB_A OUT VB_A
+ OUT OUT m9m10 OUT VCC OUT VCC VCC m9m10 m9m10 VCC m9m10 m9m10 m9m10 VB_A VB_A VB_A
+ VCC OUT VB_A VCC VB_A OUT VCC VB_A OUT VCC VB_A OUT m9m10 m9m10 m9m10 VSS sky130_fd_pr__pfet_01v8_UDM5A5
XXM9_dummy_1 dummy_9 dummy_9 bias1 VCC bias1 dummy_9 dummy_9 bias1 VCC VCC dummy_9
+ bias1 dummy_9 VCC VCC dummy_9 dummy_9 dummy_9 bias1 bias1 VCC VCC dummy_9 bias1
+ dummy_9 dummy_9 dummy_9 dummy_9 bias1 VCC dummy_9 dummy_9 bias1 VCC dummy_9 dummy_9
+ dummy_9 dummy_9 VCC bias1 VCC bias1 dummy_9 bias1 dummy_9 dummy_9 dummy_9 bias1
+ dummy_9 dummy_9 bias1 dummy_9 bias1 VCC VCC dummy_9 VCC VCC bias1 dummy_9 dummy_9
+ bias1 dummy_9 dummy_9 bias1 bias1 VCC VCC dummy_9 dummy_9 bias1 dummy_9 bias1 dummy_9
+ dummy_9 dummy_9 bias1 dummy_9 VCC VCC dummy_9 VCC VCC dummy_9 VCC dummy_9 bias1
+ dummy_9 bias1 dummy_9 bias1 bias1 bias1 VCC dummy_9 VCC bias1 dummy_9 dummy_9 dummy_9
+ dummy_9 bias1 dummy_9 dummy_9 VCC bias1 VCC VCC dummy_9 dummy_9 dummy_9 bias1 dummy_9
+ dummy_9 dummy_9 bias1 VCC bias1 dummy_9 VCC dummy_9 dummy_9 dummy_9 VCC bias1 VCC
+ dummy_9 dummy_9 dummy_9 bias1 bias1 dummy_9 dummy_9 dummy_9 dummy_9 VCC bias1 dummy_9
+ VCC dummy_9 bias1 VCC dummy_9 VCC dummy_9 dummy_9 dummy_9 VCC VCC dummy_9 VCC VCC
+ bias1 bias1 dummy_9 dummy_9 dummy_9 dummy_9 dummy_9 dummy_9 dummy_9 VCC VCC dummy_9
+ dummy_9 bias1 dummy_9 dummy_9 bias1 VCC dummy_9 dummy_9 dummy_9 dummy_9 VCC dummy_9
+ dummy_9 dummy_9 VCC VCC dummy_9 bias1 dummy_9 bias1 bias1 dummy_9 bias1 VCC dummy_9
+ bias1 VCC bias1 VCC dummy_9 VCC dummy_9 dummy_9 bias1 bias1 dummy_9 bias1 bias1
+ VCC bias1 dummy_9 dummy_9 dummy_9 VCC bias1 bias1 VCC VCC dummy_9 dummy_9 bias1
+ dummy_9 bias1 dummy_9 dummy_9 VCC bias1 dummy_9 bias1 dummy_9 dummy_9 bias1 dummy_9
+ bias1 VCC dummy_9 dummy_9 dummy_9 bias1 dummy_9 dummy_9 dummy_9 bias1 bias1 dummy_9
+ dummy_9 bias1 VCC dummy_9 dummy_9 bias1 VCC VCC dummy_9 bias1 dummy_9 bias1 dummy_9
+ bias1 VCC dummy_9 bias1 VCC dummy_9 dummy_9 bias1 dummy_9 bias1 dummy_9 dummy_9
+ VCC VCC VCC dummy_9 bias1 VCC VCC VCC dummy_9 dummy_9 dummy_9 bias1 bias1 dummy_9
+ dummy_9 VCC VCC VCC bias1 bias1 dummy_9 dummy_9 VCC VCC dummy_9 dummy_9 dummy_9
+ VCC VCC VCC VCC bias1 VCC VCC dummy_9 bias1 dummy_9 dummy_9 dummy_9 bias1 bias1
+ dummy_9 dummy_9 dummy_9 dummy_9 bias1 dummy_9 VCC VCC dummy_9 bias1 dummy_9 dummy_9
+ bias1 dummy_9 dummy_9 VCC VCC dummy_9 dummy_9 VCC dummy_9 dummy_9 bias1 dummy_9
+ dummy_9 bias1 dummy_9 dummy_9 bias1 dummy_9 VCC bias1 dummy_9 bias1 VCC dummy_9
+ bias1 VCC dummy_9 dummy_9 dummy_9 VCC VCC dummy_9 bias1 VCC dummy_9 dummy_9 bias1
+ dummy_9 VCC dummy_9 dummy_9 dummy_9 VCC bias1 dummy_9 dummy_9 VCC VCC dummy_9 bias1
+ dummy_9 bias1 dummy_9 dummy_9 dummy_9 dummy_9 dummy_9 VCC VCC dummy_9 bias1 dummy_9
+ bias1 bias1 dummy_9 bias1 dummy_9 dummy_9 VCC VCC VCC dummy_9 dummy_9 dummy_9 bias1
+ dummy_9 dummy_9 dummy_9 bias1 VCC VCC bias1 dummy_9 dummy_9 dummy_9 VCC dummy_9
+ VCC VCC VSS dummy_9 dummy_9 sky130_fd_pr__pfet_01v8_E769TZ
XXM2_dummy_9 VB_A dummy_2 VCC dummy_2 VSS sky130_fd_pr__pfet_01v8_SKU9VM
XXM5_dummy_1 VCC IN_P IN_P dummy_5 IN_P VCC dummy_5 VCC dummy_5 dummy_5 dummy_5 dummy_5
+ IN_P dummy_5 dummy_5 VCC dummy_5 IN_P dummy_5 dummy_5 VCC dummy_5 IN_P IN_P dummy_5
+ VCC IN_P IN_P IN_P VCC VCC dummy_5 VCC IN_P IN_P VCC IN_P dummy_5 dummy_5 dummy_5
+ dummy_5 IN_P VCC dummy_5 dummy_5 dummy_5 dummy_5 IN_P VCC dummy_5 dummy_5 VCC dummy_5
+ dummy_5 VCC VCC dummy_5 dummy_5 dummy_5 dummy_5 dummy_5 dummy_5 dummy_5 VCC IN_P
+ dummy_5 IN_P VCC VSS sky130_fd_pr__pfet_01v8_8DHNHY
XXM9_dummy_3 VCC bias1 dummy_9 dummy_9 VSS sky130_fd_pr__pfet_01v8_SLZ774
XXM5_dummy_3 dummy_5 IN_P VCC dummy_5 VSS sky130_fd_pr__pfet_01v8_MGA63L
XXM9_dummy_4 VCC bias1 dummy_9 dummy_9 VSS sky130_fd_pr__pfet_01v8_ZLZ7XS
XXM5_dummy_4 dummy_5 IN_P VCC dummy_5 VSS sky130_fd_pr__pfet_01v8_MGA63L
Xsky130_fd_pr__pfet_01v8_UDMRD5_0 dummy_2 dummy_2 VB_A VB_A dummy_2 dummy_2 VB_A dummy_2
+ VCC VCC dummy_2 dummy_2 dummy_2 VB_A VCC dummy_2 dummy_2 VCC dummy_2 VCC VCC VB_A
+ dummy_2 VCC VB_A dummy_2 VCC dummy_2 VB_A VB_A dummy_2 VB_A dummy_2 dummy_2 dummy_2
+ dummy_2 dummy_2 VCC dummy_2 VCC VCC dummy_2 dummy_2 VCC dummy_2 dummy_2 dummy_2
+ VB_A VB_A VB_A VCC dummy_2 VB_A VB_A VCC VB_A dummy_2 VCC VB_A dummy_2 VCC dummy_2
+ VB_A dummy_2 dummy_2 VCC dummy_2 dummy_2 VSS sky130_fd_pr__pfet_01v8_UDMRD5
XXM9_dummy_5 VCC bias1 dummy_9 dummy_9 VSS sky130_fd_pr__pfet_01v8_ZLZ7XS
XXM9_1 VCC VCC bias1 VCC bias1 VCC m9m10 bias1 VCC VCC m9m10 bias1 VCC VCC m9m10 VCC
+ m9m10 bias1 bias1 VCC VCC m9m10 bias1 VCC VCC VCC VCC bias1 VCC VCC m9m10 bias1
+ VCC m9m10 m9m10 VCC VCC VCC bias1 VCC bias1 VCC bias1 m9m10 VCC m9m10 bias1 VCC
+ m9m10 bias1 VCC VCC VCC m9m10 VCC VCC bias1 m9m10 m9m10 bias1 VCC VCC bias1 bias1
+ VCC VCC m9m10 VCC bias1 m9m10 bias1 m9m10 VCC m9m10 bias1 VCC VCC VCC m9m10 VCC
+ VCC VCC VCC VCC bias1 VCC bias1 m9m10 bias1 bias1 bias1 VCC m9m10 VCC bias1 VCC
+ m9m10 VCC m9m10 bias1 VCC VCC VCC VCC bias1 VCC VCC VCC m9m10 bias1 m9m10 VCC VCC
+ bias1 VCC bias1 m9m10 VCC VCC VCC VCC bias1 VCC m9m10 VCC m9m10 bias1 bias1 m9m10
+ m9m10 VCC VCC bias1 VCC VCC VCC bias1 VCC m9m10 m9m10 VCC VCC VCC VCC m9m10 VCC
+ VCC bias1 bias1 VCC VCC m9m10 VCC m9m10 m9m10 VCC VCC VCC m9m10 bias1 m9m10 VCC
+ bias1 VCC m9m10 VCC VCC VCC VCC m9m10 VCC m9m10 VCC VCC VCC bias1 VCC bias1 bias1
+ m9m10 bias1 VCC m9m10 bias1 VCC bias1 VCC VCC VCC VCC VCC bias1 bias1 m9m10 bias1
+ bias1 VCC bias1 m9m10 VCC VCC VCC bias1 bias1 VCC VCC VCC VCC bias1 m9m10 bias1
+ m9m10 m9m10 VCC m9m10 bias1 VCC VCC bias1 VCC bias1 VCC m9m10 m9m10 m9m10 bias1
+ VCC VCC m9m10 bias1 bias1 m9m10 m9m10 bias1 VCC m9m10 VCC bias1 VCC VCC m9m10 bias1
+ VCC bias1 m9m10 bias1 VCC m9m10 bias1 VCC m9m10 m9m10 bias1 m9m10 bias1 VCC VCC
+ VCC VCC VCC m9m10 bias1 VCC VCC VCC m9m10 m9m10 VCC bias1 bias1 m9m10 VCC VCC VCC
+ VCC bias1 bias1 m9m10 m9m10 VCC VCC VCC VCC VCC VCC VCC VCC VCC bias1 VCC VCC VCC
+ bias1 m9m10 m9m10 m9m10 bias1 bias1 m9m10 m9m10 VCC VCC bias1 VCC VCC VCC bias1
+ VCC m9m10 bias1 VCC VCC VCC VCC VCC m9m10 VCC VCC m9m10 bias1 VCC VCC bias1 VCC
+ m9m10 bias1 m9m10 VCC bias1 m9m10 bias1 VCC m9m10 bias1 VCC m9m10 m9m10 VCC VCC
+ VCC m9m10 bias1 VCC VCC m9m10 bias1 VCC VCC VCC VCC VCC VCC bias1 VCC m9m10 VCC
+ VCC m9m10 bias1 m9m10 bias1 VCC m9m10 VCC m9m10 VCC VCC VCC m9m10 bias1 m9m10 bias1
+ bias1 VCC bias1 m9m10 m9m10 VCC VCC VCC m9m10 m9m10 m9m10 bias1 m9m10 m9m10 VCC
+ bias1 VCC VCC bias1 m9m10 VCC VCC VCC VCC VCC VCC VSS m9m10 VCC sky130_fd_pr__pfet_01v8_F76D73
XXM9_dummy_20 VCC bias1 dummy_9 dummy_9 VSS sky130_fd_pr__pfet_01v8_ZLZ7XS
XXM5_dummy_5 dummy_5 IN_P VCC dummy_5 VSS sky130_fd_pr__pfet_01v8_MGA63L
XXM9_dummy_6 VCC bias1 dummy_9 dummy_9 VSS sky130_fd_pr__pfet_01v8_ZLZ7XS
XXM9_dummy_10 VCC bias1 dummy_9 dummy_9 VSS sky130_fd_pr__pfet_01v8_ZLZ7XS
XXM9_2 VCC VCC bias1 VCC bias1 VCC m9m10 bias1 VCC VCC m9m10 bias1 VCC VCC m9m10 VCC
+ m9m10 bias1 bias1 VCC VCC m9m10 bias1 VCC VCC VCC VCC bias1 VCC VCC m9m10 bias1
+ VCC m9m10 m9m10 VCC VCC VCC bias1 VCC bias1 VCC bias1 m9m10 VCC m9m10 bias1 VCC
+ m9m10 bias1 VCC VCC VCC m9m10 VCC VCC bias1 m9m10 m9m10 bias1 VCC VCC bias1 bias1
+ VCC VCC m9m10 VCC bias1 m9m10 bias1 m9m10 VCC m9m10 bias1 VCC VCC VCC m9m10 VCC
+ VCC VCC VCC VCC bias1 VCC bias1 m9m10 bias1 bias1 bias1 VCC m9m10 VCC bias1 VCC
+ m9m10 VCC m9m10 bias1 VCC VCC VCC VCC bias1 VCC VCC VCC m9m10 bias1 m9m10 VCC VCC
+ bias1 VCC bias1 m9m10 VCC VCC VCC VCC bias1 VCC m9m10 VCC m9m10 bias1 bias1 m9m10
+ m9m10 VCC VCC bias1 VCC VCC VCC bias1 VCC m9m10 m9m10 VCC VCC VCC VCC m9m10 VCC
+ VCC bias1 bias1 VCC VCC m9m10 VCC m9m10 m9m10 VCC VCC VCC m9m10 bias1 m9m10 VCC
+ bias1 VCC m9m10 VCC VCC VCC VCC m9m10 VCC m9m10 VCC VCC VCC bias1 VCC bias1 bias1
+ m9m10 bias1 VCC m9m10 bias1 VCC bias1 VCC VCC VCC VCC VCC bias1 bias1 m9m10 bias1
+ bias1 VCC bias1 m9m10 VCC VCC VCC bias1 bias1 VCC VCC VCC VCC bias1 m9m10 bias1
+ m9m10 m9m10 VCC m9m10 bias1 VCC VCC bias1 VCC bias1 VCC m9m10 m9m10 m9m10 bias1
+ VCC VCC m9m10 bias1 bias1 m9m10 m9m10 bias1 VCC m9m10 VCC bias1 VCC VCC m9m10 bias1
+ VCC bias1 m9m10 bias1 VCC m9m10 bias1 VCC m9m10 m9m10 bias1 m9m10 bias1 VCC VCC
+ VCC VCC VCC m9m10 bias1 VCC VCC VCC m9m10 m9m10 VCC bias1 bias1 m9m10 VCC VCC VCC
+ VCC bias1 bias1 m9m10 m9m10 VCC VCC VCC VCC VCC VCC VCC VCC VCC bias1 VCC VCC VCC
+ bias1 m9m10 m9m10 m9m10 bias1 bias1 m9m10 m9m10 VCC VCC bias1 VCC VCC VCC bias1
+ VCC m9m10 bias1 VCC VCC VCC VCC VCC m9m10 VCC VCC m9m10 bias1 VCC VCC bias1 VCC
+ m9m10 bias1 m9m10 VCC bias1 m9m10 bias1 VCC m9m10 bias1 VCC m9m10 m9m10 VCC VCC
+ VCC m9m10 bias1 VCC VCC m9m10 bias1 VCC VCC VCC VCC VCC VCC bias1 VCC m9m10 VCC
+ VCC m9m10 bias1 m9m10 bias1 VCC m9m10 VCC m9m10 VCC VCC VCC m9m10 bias1 m9m10 bias1
+ bias1 VCC bias1 m9m10 m9m10 VCC VCC VCC m9m10 m9m10 m9m10 bias1 m9m10 m9m10 VCC
+ bias1 VCC VCC bias1 m9m10 VCC VCC VCC VCC VCC VCC VSS m9m10 VCC sky130_fd_pr__pfet_01v8_F76D73
XXM5_dummy_6 dummy_5 IN_P VCC dummy_5 VSS sky130_fd_pr__pfet_01v8_MGA63L
XXM9_dummy_7 VCC bias1 dummy_9 dummy_9 VSS sky130_fd_pr__pfet_01v8_ZLZ7XS
XXM9_dummy_22 VCC bias1 dummy_9 dummy_9 VSS sky130_fd_pr__pfet_01v8_ZLZ7XS
XXM9_dummy_11 VCC bias1 dummy_9 dummy_9 VSS sky130_fd_pr__pfet_01v8_ZLZ7XS
XXM9_3 VCC VCC bias1 VCC bias1 VCC m9m10 bias1 VCC VCC m9m10 bias1 VCC VCC m9m10 VCC
+ m9m10 bias1 bias1 VCC VCC m9m10 bias1 VCC VCC VCC VCC bias1 VCC VCC m9m10 bias1
+ VCC m9m10 m9m10 VCC VCC VCC bias1 VCC bias1 VCC bias1 m9m10 VCC m9m10 bias1 VCC
+ m9m10 bias1 VCC VCC VCC m9m10 VCC VCC bias1 m9m10 m9m10 bias1 VCC VCC bias1 bias1
+ VCC VCC m9m10 VCC bias1 m9m10 bias1 m9m10 VCC m9m10 bias1 VCC VCC VCC m9m10 VCC
+ VCC VCC VCC VCC bias1 VCC bias1 m9m10 bias1 bias1 bias1 VCC m9m10 VCC bias1 VCC
+ m9m10 VCC m9m10 bias1 VCC VCC VCC VCC bias1 VCC VCC VCC m9m10 bias1 m9m10 VCC VCC
+ bias1 VCC bias1 m9m10 VCC VCC VCC VCC bias1 VCC m9m10 VCC m9m10 bias1 bias1 m9m10
+ m9m10 VCC VCC bias1 VCC VCC VCC bias1 VCC m9m10 m9m10 VCC VCC VCC VCC m9m10 VCC
+ VCC bias1 bias1 VCC VCC m9m10 VCC m9m10 m9m10 VCC VCC VCC m9m10 bias1 m9m10 VCC
+ bias1 VCC m9m10 VCC VCC VCC VCC m9m10 VCC m9m10 VCC VCC VCC bias1 VCC bias1 bias1
+ m9m10 bias1 VCC m9m10 bias1 VCC bias1 VCC VCC VCC VCC VCC bias1 bias1 m9m10 bias1
+ bias1 VCC bias1 m9m10 VCC VCC VCC bias1 bias1 VCC VCC VCC VCC bias1 m9m10 bias1
+ m9m10 m9m10 VCC m9m10 bias1 VCC VCC bias1 VCC bias1 VCC m9m10 m9m10 m9m10 bias1
+ VCC VCC m9m10 bias1 bias1 m9m10 m9m10 bias1 VCC m9m10 VCC bias1 VCC VCC m9m10 bias1
+ VCC bias1 m9m10 bias1 VCC m9m10 bias1 VCC m9m10 m9m10 bias1 m9m10 bias1 VCC VCC
+ VCC VCC VCC m9m10 bias1 VCC VCC VCC m9m10 m9m10 VCC bias1 bias1 m9m10 VCC VCC VCC
+ VCC bias1 bias1 m9m10 m9m10 VCC VCC VCC VCC VCC VCC VCC VCC VCC bias1 VCC VCC VCC
+ bias1 m9m10 m9m10 m9m10 bias1 bias1 m9m10 m9m10 VCC VCC bias1 VCC VCC VCC bias1
+ VCC m9m10 bias1 VCC VCC VCC VCC VCC m9m10 VCC VCC m9m10 bias1 VCC VCC bias1 VCC
+ m9m10 bias1 m9m10 VCC bias1 m9m10 bias1 VCC m9m10 bias1 VCC m9m10 m9m10 VCC VCC
+ VCC m9m10 bias1 VCC VCC m9m10 bias1 VCC VCC VCC VCC VCC VCC bias1 VCC m9m10 VCC
+ VCC m9m10 bias1 m9m10 bias1 VCC m9m10 VCC m9m10 VCC VCC VCC m9m10 bias1 m9m10 bias1
+ bias1 VCC bias1 m9m10 m9m10 VCC VCC VCC m9m10 m9m10 m9m10 bias1 m9m10 m9m10 VCC
+ bias1 VCC VCC bias1 m9m10 VCC VCC VCC VCC VCC VCC VSS m9m10 VCC sky130_fd_pr__pfet_01v8_F76D73
XXM11_1 OUT OUT VB_B OUT VB_B VB_B VB_B VB_B m11m12 m11m12 m11m12 m11m12 OUT OUT VB_B
+ OUT OUT VB_B OUT OUT m11m12 VB_B m11m12 m11m12 m11m12 m11m12 m11m12 VB_B VB_B OUT
+ OUT VB_B OUT VB_B OUT VB_B VB_B m11m12 VB_B m11m12 m11m12 m11m12 m11m12 OUT OUT
+ VSS sky130_fd_pr__nfet_01v8_QP5WRD
XXM5_dummy_7 dummy_5 IN_P VCC dummy_5 VSS sky130_fd_pr__pfet_01v8_MGA63L
XXM9_dummy_8 VCC bias1 dummy_9 dummy_9 VSS sky130_fd_pr__pfet_01v8_ZLZ7XS
Xsky130_fd_pr__nfet_01v8_SCE452_0 dummy_4 bias3 dummy_4 VSS sky130_fd_pr__nfet_01v8_SCE452
XXM9_4 VCC VCC bias1 VCC bias1 VCC m9m10 bias1 VCC VCC m9m10 bias1 VCC VCC m9m10 VCC
+ m9m10 bias1 bias1 VCC VCC m9m10 bias1 VCC VCC VCC VCC bias1 VCC VCC m9m10 bias1
+ VCC m9m10 m9m10 VCC VCC VCC bias1 VCC bias1 VCC bias1 m9m10 VCC m9m10 bias1 VCC
+ m9m10 bias1 VCC VCC VCC m9m10 VCC VCC bias1 m9m10 m9m10 bias1 VCC VCC bias1 bias1
+ VCC VCC m9m10 VCC bias1 m9m10 bias1 m9m10 VCC m9m10 bias1 VCC VCC VCC m9m10 VCC
+ VCC VCC VCC VCC bias1 VCC bias1 m9m10 bias1 bias1 bias1 VCC m9m10 VCC bias1 VCC
+ m9m10 VCC m9m10 bias1 VCC VCC VCC VCC bias1 VCC VCC VCC m9m10 bias1 m9m10 VCC VCC
+ bias1 VCC bias1 m9m10 VCC VCC VCC VCC bias1 VCC m9m10 VCC m9m10 bias1 bias1 m9m10
+ m9m10 VCC VCC bias1 VCC VCC VCC bias1 VCC m9m10 m9m10 VCC VCC VCC VCC m9m10 VCC
+ VCC bias1 bias1 VCC VCC m9m10 VCC m9m10 m9m10 VCC VCC VCC m9m10 bias1 m9m10 VCC
+ bias1 VCC m9m10 VCC VCC VCC VCC m9m10 VCC m9m10 VCC VCC VCC bias1 VCC bias1 bias1
+ m9m10 bias1 VCC m9m10 bias1 VCC bias1 VCC VCC VCC VCC VCC bias1 bias1 m9m10 bias1
+ bias1 VCC bias1 m9m10 VCC VCC VCC bias1 bias1 VCC VCC VCC VCC bias1 m9m10 bias1
+ m9m10 m9m10 VCC m9m10 bias1 VCC VCC bias1 VCC bias1 VCC m9m10 m9m10 m9m10 bias1
+ VCC VCC m9m10 bias1 bias1 m9m10 m9m10 bias1 VCC m9m10 VCC bias1 VCC VCC m9m10 bias1
+ VCC bias1 m9m10 bias1 VCC m9m10 bias1 VCC m9m10 m9m10 bias1 m9m10 bias1 VCC VCC
+ VCC VCC VCC m9m10 bias1 VCC VCC VCC m9m10 m9m10 VCC bias1 bias1 m9m10 VCC VCC VCC
+ VCC bias1 bias1 m9m10 m9m10 VCC VCC VCC VCC VCC VCC VCC VCC VCC bias1 VCC VCC VCC
+ bias1 m9m10 m9m10 m9m10 bias1 bias1 m9m10 m9m10 VCC VCC bias1 VCC VCC VCC bias1
+ VCC m9m10 bias1 VCC VCC VCC VCC VCC m9m10 VCC VCC m9m10 bias1 VCC VCC bias1 VCC
+ m9m10 bias1 m9m10 VCC bias1 m9m10 bias1 VCC m9m10 bias1 VCC m9m10 m9m10 VCC VCC
+ VCC m9m10 bias1 VCC VCC m9m10 bias1 VCC VCC VCC VCC VCC VCC bias1 VCC m9m10 VCC
+ VCC m9m10 bias1 m9m10 bias1 VCC m9m10 VCC m9m10 VCC VCC VCC m9m10 bias1 m9m10 bias1
+ bias1 VCC bias1 m9m10 m9m10 VCC VCC VCC m9m10 m9m10 m9m10 bias1 m9m10 m9m10 VCC
+ bias1 VCC VCC bias1 m9m10 VCC VCC VCC VCC VCC VCC VSS m9m10 VCC sky130_fd_pr__pfet_01v8_F76D73
XXM9_dummy_12 VCC bias1 dummy_9 dummy_9 VSS sky130_fd_pr__pfet_01v8_ZLZ7XS
XXM5_dummy_8 dummy_5 IN_P VCC dummy_5 VSS sky130_fd_pr__pfet_01v8_MGA63L
XXM9_dummy_9 VCC bias1 dummy_9 dummy_9 VSS sky130_fd_pr__pfet_01v8_ZLZ7XS
XXM10 OUT VB_A m9m10 OUT VB_A m9m10 VCC VCC m9m10 m9m10 m9m10 VB_A VCC m9m10 VCC OUT
+ VCC VCC VB_A OUT VCC VB_A OUT OUT VB_A VB_A m9m10 VB_A m9m10 m9m10 OUT m9m10 VCC
+ m9m10 VCC VCC OUT OUT VCC OUT OUT OUT VB_A VB_A VB_A VCC m9m10 VB_A VCC VB_A m9m10
+ VCC VB_A m9m10 VCC VB_A m9m10 OUT OUT OUT VSS sky130_fd_pr__pfet_01v8_UDM5A5
Xsky130_fd_pr__nfet_01v8_SCE452_1 dummy_4 bias3 dummy_4 VSS sky130_fd_pr__nfet_01v8_SCE452
Xsky130_fd_pr__pfet_01v8_7DHACV_0 VCC IN_P IN_P m1_44990_37960# VCC VCC bias21 bias21
+ bias21 m1_44990_37960# IN_P m1_44990_37960# bias21 m1_44990_37960# IN_P bias21 m1_44990_37960#
+ VCC IN_P IN_P m1_44990_37960# VCC IN_P IN_P IN_P VCC VCC VCC IN_P IN_P IN_P bias21
+ bias21 bias21 m1_44990_37960# IN_P VCC m1_44990_37960# bias21 m1_44990_37960# bias21
+ IN_P VCC m1_44990_37960# bias21 VCC m1_44990_37960# VCC VCC bias21 m1_44990_37960#
+ bias21 m1_44990_37960# m1_44990_37960# bias21 m1_44990_37960# VCC bias21 IN_P VCC
+ VSS sky130_fd_pr__pfet_01v8_7DHACV
XXM9_dummy_13 VCC bias1 dummy_9 dummy_9 VSS sky130_fd_pr__pfet_01v8_ZLZ7XS
XXM100_1 IB VCC VCC m1_44990_37960# VCC IB m1_44990_37960# IB VCC m1_44990_37960#
+ VCC VCC VSS sky130_fd_pr__pfet_01v8_RRU5GE
XXM2_dummy_10 VB_A dummy_2 VCC dummy_2 VSS sky130_fd_pr__pfet_01v8_SKU9VM
XXM11 m11m12 m11m12 VB_B m11m12 VB_B VB_B VB_B VB_B OUT OUT OUT OUT m11m12 m11m12
+ VB_B m11m12 m11m12 VB_B m11m12 m11m12 OUT VB_B OUT OUT OUT OUT OUT VB_B VB_B m11m12
+ m11m12 VB_B m11m12 VB_B m11m12 VB_B VB_B OUT VB_B OUT OUT OUT OUT m11m12 m11m12
+ VSS sky130_fd_pr__nfet_01v8_QP5WRD
Xsky130_fd_pr__nfet_01v8_SCE452_2 dummy_4 bias3 dummy_4 VSS sky130_fd_pr__nfet_01v8_SCE452
Xsky130_fd_pr__nfet_01v8_WK8VRD_0 VB_B dummy_3 dummy_3 dummy_3 VB_B dummy_3 VB_B VB_B
+ VB_B VB_B dummy_3 dummy_3 dummy_3 dummy_3 dummy_3 dummy_3 VB_B dummy_3 dummy_3 dummy_3
+ VB_B dummy_3 dummy_3 dummy_3 VB_B dummy_3 dummy_3 dummy_3 dummy_3 VB_B dummy_3 dummy_3
+ VB_B VB_B dummy_3 dummy_3 VB_B dummy_3 VB_B dummy_3 VB_B VB_B dummy_3 VB_B dummy_3
+ dummy_3 dummy_3 dummy_3 dummy_3 dummy_3 dummy_3 VSS sky130_fd_pr__nfet_01v8_WK8VRD
XXM9_dummy_14 VCC bias1 dummy_9 dummy_9 VSS sky130_fd_pr__pfet_01v8_ZLZ7XS
C0 dummy_5 VCC 11.5f
C1 VB_A dummy_2 33f
C2 dummy_4 m11m12 1.08f
C3 bias21 dummy_4 0.403f
C4 m11m12 bias3 0.374f
C5 VB_A bias1 7.09f
C6 bias21 bias3 10.1f
C7 VB_B m3m4 6.64f
C8 IN_P m1_44990_37960# 13.5f
C9 dummy_2 VCC 13f
C10 m1m2 VB_A 6.26f
C11 OUT bias3 0.978f
C12 VCC bias1 0.898p
C13 dummy_5 bias3 0.399f
C14 bias21 m11m12 0.836f
C15 m1m2 VCC 0.153p
C16 OUT m11m12 -1.26f
C17 dummy_3 m11m12 20.7f
C18 bias1 dummy_9 0.104p
C19 OUT bias21 0.978f
C20 IB VCC 25.7f
C21 IN_M m1_44990_37960# 10.4f
C22 dummy_3 bias21 0.965f
C23 dummy_100 VCC 8.42f
C24 m1m2 dummy_9 35f
C25 OUT dummy_3 2.64f
C26 dummy_5 bias21 0.398f
C27 m1_44990_37960# VCC 31.6f
C28 VB_A m9m10 5.59f
C29 bias21 dummy_2 0.891f
C30 m9m10 VCC 0.147p
C31 OUT dummy_2 15.7f
C32 IN_P IN_M 3.48f
C33 IB bias3 0.799f
C34 VB_B VCC 2.87f
C35 m9m10 dummy_9 35.9f
C36 dummy_4 m3m4 1.44f
C37 IN_P VCC 29.4f
C38 m1_44990_37960# bias3 0.988f
C39 OUT bias1 1.55f
C40 dummy_3 bias1 2.66f
C41 m1m2 OUT 0.00992f
C42 bias3 m3m4 1.29f
C43 bias21 IB 0.799f
C44 bias21 m1_44990_37960# 1.69f
C45 VB_A VCC 33.9f
C46 IN_M VCC 12.3f
C47 m11m12 m3m4 0.403f
C48 VB_B bias3 0.978f
C49 bias21 m3m4 0.0154f
C50 dummy_2 bias1 2.5f
C51 OUT m3m4 18.9f
C52 dummy_3 m3m4 2.84f
C53 IN_P bias3 0.727f
C54 dummy_5 m1_44990_37960# 15.6f
C55 m1m2 dummy_2 2.66f
C56 VB_B m11m12 6.51f
C57 VB_B bias21 1.01f
C58 OUT m9m10 -1.25f
C59 VCC dummy_9 0.127p
C60 m1m2 bias1 61.6f
C61 OUT VB_B 5.56f
C62 VB_B dummy_3 33.2f
C63 IN_P bias21 11.1f
C64 VB_A bias3 0.978f
C65 IN_M bias3 10.4f
C66 IN_P dummy_5 31.3f
C67 dummy_100 IB 16.7f
C68 bias3 VCC 41.2f
C69 bias21 VB_A 1.01f
C70 m3m4 bias1 -1.25f
C71 dummy_2 m9m10 2.69f
C72 OUT VB_A 6.54f
C73 IB m1_44990_37960# 7.64f
C74 dummy_100 m1_44990_37960# 5.9f
C75 m9m10 bias1 81.2f
C76 bias21 VCC 39.6f
C77 VB_B bias1 5.61f
C78 dummy_5 IN_M 2.85f
C79 OUT VCC 12.4f
C80 m1m2 m9m10 0.118p
C81 dummy_4 bias3 8.54f
C82 dummy_4 VSS 3.54f
C83 bias21 VSS 1.61f
C84 OUT VSS 26.9f
C85 m11m12 VSS 24.7f
C86 VCC VSS 22.5p
C87 dummy_5 VSS 17.1f
C88 IN_P VSS 12.5f
C89 dummy_9 VSS 0.175p
C90 bias1 VSS 3.55p
C91 m9m10 VSS 0.169p
C92 dummy_2 VSS 25.9f
C93 VB_A VSS 0.102p
C94 bias3 VSS 48.6f
C95 m1_44990_37960# VSS 8.85f
C96 IN_M VSS 8.73f
C97 m3m4 VSS 19.8f
C98 m1m2 VSS 0.157p
C99 dummy_3 VSS 43.3f
C100 VB_B VSS 0.189p
C101 dummy_100 VSS 8.79f
C102 IB VSS 25.4f
.ends

