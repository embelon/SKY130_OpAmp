VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS

LAYER via2
  TYPE CUT ;
END via2

LAYER via
  TYPE CUT ;
END via

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER via3
  TYPE CUT ;
END via3

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER via4
  TYPE CUT ;
END via4

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met6
  TYPE ROUTING ;
END met6

LAYER met1
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  DIRECTION HORIZONTAL ;
END met1

LAYER met3
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  DIRECTION HORIZONTAL ;
END met3

LAYER met2
  TYPE ROUTING ;
  WIDTH 0.140000 ;
  DIRECTION HORIZONTAL ;
END met2

LAYER met4
  TYPE ROUTING ;
  WIDTH 0.300000 ;
  DIRECTION HORIZONTAL ;
END met4

LAYER met5
  TYPE ROUTING ;
  WIDTH 1.600000 ;
  DIRECTION HORIZONTAL ;
END met5

LAYER li1
  TYPE ROUTING ;
  WIDTH 0.170000 ;
  DIRECTION HORIZONTAL ;
END li1

MACRO opamp_cascode
  CLASS BLOCK ;
  FOREIGN opamp_cascode ;
  ORIGIN -170.000 -70.000 ;
  SIZE 360.000 BY 650.000 ;
  PIN IN_P
    ANTENNAGATEAREA 64.799995 ;
    PORT
      LAYER met2 ;
        RECT 170.000 71.000 171.000 80.000 ;
        RECT 170.000 70.000 180.000 71.000 ;
    END
  END IN_P
  PIN IN_M
    ANTENNAGATEAREA 27.000000 ;
    PORT
      LAYER met2 ;
        RECT 170.000 90.000 171.000 100.000 ;
    END
  END IN_M
  PIN VCC
    ANTENNADIFFAREA 1468.099976 ;
    PORT
      LAYER nwell ;
        RECT 300.000 719.000 530.000 720.000 ;
        RECT 170.000 430.000 171.000 440.000 ;
        RECT 170.000 270.000 171.000 280.000 ;
        RECT 529.000 71.000 530.000 719.000 ;
        RECT 190.000 70.000 530.000 71.000 ;
      LAYER met2 ;
        RECT 170.000 719.000 180.000 720.000 ;
        RECT 170.000 710.000 171.000 719.000 ;
    END
  END VCC
  PIN VSS
    ANTENNADIFFAREA 21.400000 ;
    PORT
      LAYER pwell ;
        RECT 190.000 719.000 284.000 720.000 ;
        RECT 170.000 560.000 171.000 570.000 ;
      LAYER met2 ;
        RECT 170.000 660.000 171.000 670.000 ;
    END
  END VSS
  PIN OUT
    ANTENNADIFFAREA 87.000000 ;
    PORT
      LAYER met2 ;
        RECT 170.000 450.000 171.000 460.000 ;
    END
  END OUT
  PIN VB_A
    ANTENNAGATEAREA 2550.000000 ;
    PORT
      LAYER met2 ;
        RECT 170.000 430.000 171.000 440.000 ;
    END
  END VB_A
  PIN VB_B
    ANTENNAGATEAREA 2550.000000 ;
    PORT
      LAYER met2 ;
        RECT 170.000 560.000 171.000 570.000 ;
    END
  END VB_B
  PIN IB
    ANTENNAGATEAREA 450.000000 ;
    ANTENNADIFFAREA 5.800000 ;
    PORT
      LAYER met2 ;
        RECT 170.000 270.000 171.000 280.000 ;
    END
  END IB
  OBS
      LAYER li1 ;
        RECT 300.700 719.000 304.300 719.400 ;
        RECT 201.500 79.095 523.700 719.000 ;
      LAYER mcon ;
        RECT 300.700 718.800 304.300 719.400 ;
      LAYER met1 ;
        RECT 170.000 719.000 490.000 720.000 ;
        RECT 170.000 710.000 524.500 719.000 ;
        RECT 171.000 670.000 524.500 710.000 ;
        RECT 170.000 660.000 524.500 670.000 ;
        RECT 171.000 570.000 524.500 660.000 ;
        RECT 170.000 560.000 524.500 570.000 ;
        RECT 171.000 460.075 524.500 560.000 ;
        RECT 170.000 450.000 524.500 460.075 ;
        RECT 171.000 440.000 524.500 450.000 ;
        RECT 170.000 430.000 524.500 440.000 ;
        RECT 171.000 280.000 524.500 430.000 ;
        RECT 170.000 270.000 524.500 280.000 ;
        RECT 171.000 100.000 524.500 270.000 ;
        RECT 170.000 90.000 524.500 100.000 ;
        RECT 171.000 80.000 524.500 90.000 ;
        RECT 170.000 71.000 524.500 80.000 ;
        RECT 170.000 70.000 180.000 71.000 ;
      LAYER met2 ;
        RECT 171.000 71.000 524.000 719.000 ;
  END
END opamp_cascode
END LIBRARY

