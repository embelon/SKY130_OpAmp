VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO opamp_cascode
  CLASS BLOCK ;
  FOREIGN opamp_cascode ;
  ORIGIN -164.000 -70.000 ;
  SIZE 366.000 BY 655.000 ;
  PIN IN_P
    ANTENNAGATEAREA 64.799995 ;
    PORT
      LAYER met3 ;
        RECT 166.800 71.600 167.800 72.600 ;
    END
  END IN_P
  PIN IN_M
    ANTENNAGATEAREA 27.000000 ;
    PORT
      LAYER met3 ;
        RECT 168.300 92.800 169.300 93.800 ;
    END
  END IN_M
  PIN VCC
    ANTENNADIFFAREA 1468.099976 ;
    PORT
      LAYER met3 ;
        RECT 167.600 699.100 168.600 700.100 ;
    END
  END VCC
  PIN VSS
    ANTENNADIFFAREA 21.400000 ;
    PORT
      LAYER met3 ;
        RECT 166.700 717.200 167.700 718.200 ;
    END
  END VSS
  PIN OUT
    ANTENNADIFFAREA 87.000000 ;
    PORT
      LAYER met3 ;
        RECT 168.025 453.320 169.025 454.320 ;
    END
  END OUT
  PIN VB_A
    ANTENNAGATEAREA 2550.000000 ;
    PORT
      LAYER met3 ;
        RECT 167.500 432.400 168.500 433.400 ;
    END
  END VB_A
  PIN VB_B
    ANTENNAGATEAREA 2550.000000 ;
    PORT
      LAYER met3 ;
        RECT 167.300 565.300 168.300 566.300 ;
    END
  END VB_B
  PIN IB
    ANTENNAGATEAREA 450.000000 ;
    ANTENNADIFFAREA 5.800000 ;
    PORT
      LAYER met3 ;
        RECT 164.700 272.200 165.700 273.200 ;
    END
  END IB
  OBS
      LAYER li1 ;
        RECT 201.500 79.095 523.700 719.400 ;
      LAYER met1 ;
        RECT 201.950 74.500 524.500 722.000 ;
      LAYER met2 ;
        RECT 180.000 71.950 524.000 725.000 ;
      LAYER met3 ;
        RECT 164.000 718.200 273.050 725.000 ;
        RECT 164.000 717.200 166.700 718.200 ;
        RECT 168.100 717.200 273.050 718.200 ;
        RECT 164.000 700.100 273.050 717.200 ;
        RECT 164.000 699.100 167.600 700.100 ;
        RECT 169.000 699.100 273.050 700.100 ;
        RECT 164.000 566.300 273.050 699.100 ;
        RECT 164.000 565.300 167.300 566.300 ;
        RECT 168.700 565.300 273.050 566.300 ;
        RECT 164.000 454.320 273.050 565.300 ;
        RECT 164.000 453.320 168.025 454.320 ;
        RECT 169.425 453.320 273.050 454.320 ;
        RECT 164.000 433.400 273.050 453.320 ;
        RECT 164.000 432.400 167.500 433.400 ;
        RECT 168.900 432.400 273.050 433.400 ;
        RECT 164.000 273.200 273.050 432.400 ;
        RECT 164.000 272.200 164.700 273.200 ;
        RECT 166.100 272.200 273.050 273.200 ;
        RECT 164.000 93.800 273.050 272.200 ;
        RECT 164.000 92.800 168.300 93.800 ;
        RECT 169.700 92.800 273.050 93.800 ;
        RECT 164.000 72.600 273.050 92.800 ;
        RECT 164.000 71.600 166.800 72.600 ;
        RECT 168.200 71.600 273.050 72.600 ;
        RECT 164.000 70.000 273.050 71.600 ;
  END
END opamp_cascode
END LIBRARY

