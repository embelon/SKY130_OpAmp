* NGSPICE file created from opamp_cascode.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_SCE452 a_n158_n125# a_n100_n213# a_100_n125# VSUBS
X0 a_100_n125# a_n100_n213# a_n158_n125# VSUBS sky130_fd_pr__nfet_01v8 ad=0.363 pd=3.08 as=0.363 ps=3.08 w=1.25 l=1
**devattr s=14500,616 d=14500,616
C0 a_n158_n125# a_100_n125# 0.0693f
C1 a_n100_n213# a_100_n125# 0.0322f
C2 a_n100_n213# a_n158_n125# 0.0322f
C3 a_100_n125# VSUBS 0.151f
C4 a_n158_n125# VSUBS 0.151f
C5 a_n100_n213# VSUBS 0.664f
.ends

.subckt sky130_fd_pr__pfet_01v8_ZLZ7XS w_n1594_n600# a_n1500_n597# a_1500_n500# a_n1558_n500#
+ VSUBS
X0 a_1500_n500# a_n1500_n597# a_n1558_n500# w_n1594_n600# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
C0 w_n1594_n600# a_1500_n500# 0.0187f
C1 a_n1500_n597# a_n1558_n500# 0.217f
C2 a_1500_n500# a_n1500_n597# 0.217f
C3 w_n1594_n600# a_n1558_n500# 0.0187f
C4 w_n1594_n600# a_n1500_n597# 1.65f
C5 a_1500_n500# VSUBS 0.65f
C6 a_n1558_n500# VSUBS 0.65f
C7 a_n1500_n597# VSUBS 6.74f
C8 w_n1594_n600# VSUBS 11.5f
.ends

.subckt sky130_fd_pr__pfet_01v8_7DHACV w_n112_636# a_n33_n5541# a_n33_n8013# a_n76_736#
+ w_n112_1872# w_n112_4344# a_18_n500# a_18_n2972# a_18_n5444# a_n76_n1736# a_n33_3111#
+ a_n76_n4208# a_18_3208# a_n76_n7916# a_n33_n1833# a_18_6916# a_n76_5680# w_n112_n3072#
+ a_n33_n4305# a_n33_5583# a_n76_8152# w_n112_n6780# a_n33_8055# a_n33_n3069# a_n33_639#
+ w_n112_n9252# w_n112_3108# w_n112_6816# a_n33_n6777# a_n33_n597# a_n33_n9249# a_18_n1736#
+ a_18_n4208# a_18_n7916# a_n76_1972# a_n33_1875# w_n112_n600# a_n76_n6680# a_18_736#
+ a_n76_4444# a_18_5680# a_n33_4347# w_n112_n5544# a_n76_n9152# a_18_8152# w_n112_n8016#
+ a_n76_n500# w_n112_5580# w_n112_8052# a_18_n6680# a_n76_n2972# a_18_1972# a_n76_3208#
+ a_n76_n5444# a_18_4444# a_n76_6916# w_n112_n1836# a_18_n9152# a_n33_6819# w_n112_n4308#
+ VSUBS
X0 a_18_3208# a_n33_3111# a_n76_3208# w_n112_3108# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X1 a_18_n6680# a_n33_n6777# a_n76_n6680# w_n112_n6780# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X2 a_18_n500# a_n33_n597# a_n76_n500# w_n112_n600# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X3 a_18_n9152# a_n33_n9249# a_n76_n9152# w_n112_n9252# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X4 a_18_736# a_n33_639# a_n76_736# w_n112_636# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X5 a_18_n2972# a_n33_n3069# a_n76_n2972# w_n112_n3072# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X6 a_18_n7916# a_n33_n8013# a_n76_n7916# w_n112_n8016# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X7 a_18_5680# a_n33_5583# a_n76_5680# w_n112_5580# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X8 a_18_n5444# a_n33_n5541# a_n76_n5444# w_n112_n5544# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X9 a_18_8152# a_n33_8055# a_n76_8152# w_n112_8052# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X10 a_18_n1736# a_n33_n1833# a_n76_n1736# w_n112_n1836# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X11 a_18_6916# a_n33_6819# a_n76_6916# w_n112_6816# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X12 a_18_1972# a_n33_1875# a_n76_1972# w_n112_1872# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X13 a_18_n4208# a_n33_n4305# a_n76_n4208# w_n112_n4308# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X14 a_18_4444# a_n33_4347# a_n76_4444# w_n112_4344# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
C0 w_n112_n5544# a_n33_n6777# 4.13e-19
C1 a_18_n4208# w_n112_n3072# 0.00199f
C2 w_n112_n4308# a_18_n4208# 0.0182f
C3 a_n33_n597# a_n76_n1736# 1.15e-19
C4 a_n33_8055# w_n112_6816# 4.13e-19
C5 a_n33_n4305# a_n76_n4208# 0.0417f
C6 a_18_4444# w_n112_4344# 0.0182f
C7 a_n33_4347# a_n33_5583# 0.0665f
C8 a_n76_n6680# a_n33_n5541# 1.15e-19
C9 w_n112_636# a_n33_639# 0.106f
C10 a_n33_5583# w_n112_4344# 4.13e-19
C11 a_n76_6916# a_n33_5583# 1.15e-19
C12 a_n76_n1736# w_n112_n1836# 0.0182f
C13 a_n33_n1833# w_n112_n3072# 4.13e-19
C14 w_n112_1872# a_n33_639# 4.13e-19
C15 a_n33_n8013# a_n76_n7916# 0.0417f
C16 w_n112_n5544# a_18_n6680# 0.00199f
C17 w_n112_n6780# a_n76_n6680# 0.0182f
C18 a_n33_4347# a_n76_3208# 1.15e-19
C19 a_n33_1875# a_n76_736# 1.15e-19
C20 a_n76_1972# a_n33_639# 1.15e-19
C21 a_n76_n4208# a_18_n4208# 0.747f
C22 a_n76_4444# a_18_4444# 0.747f
C23 a_n33_4347# a_n33_3111# 0.0665f
C24 a_n76_n500# a_n76_n1736# 0.00947f
C25 w_n112_n4308# a_n33_n5541# 4.13e-19
C26 a_n76_8152# w_n112_6816# 0.00199f
C27 a_18_736# a_n33_n597# 1.15e-19
C28 w_n112_n8016# a_n76_n7916# 0.0182f
C29 w_n112_n9252# a_n33_n8013# 4.13e-19
C30 a_n76_3208# w_n112_4344# 0.00199f
C31 a_18_8152# a_18_6916# 0.00947f
C32 a_n33_3111# w_n112_4344# 4.13e-19
C33 a_n76_4444# a_n33_5583# 1.15e-19
C34 a_n76_n5444# a_n76_n6680# 0.00947f
C35 a_18_n5444# a_n33_n6777# 1.15e-19
C36 a_18_n1736# w_n112_n3072# 0.00199f
C37 w_n112_n5544# a_n33_n4305# 4.13e-19
C38 w_n112_636# a_n76_736# 0.0182f
C39 a_n76_n7916# a_18_n7916# 0.747f
C40 a_n33_639# w_n112_n600# 4.13e-19
C41 a_18_6916# a_n33_5583# 1.15e-19
C42 w_n112_1872# a_n76_736# 0.00199f
C43 a_n33_6819# w_n112_8052# 4.13e-19
C44 w_n112_n4308# a_n76_n5444# 0.00199f
C45 w_n112_n9252# a_18_n7916# 0.00199f
C46 a_n76_4444# a_n76_3208# 0.00947f
C47 a_n33_4347# a_18_3208# 1.15e-19
C48 a_n76_1972# a_n76_736# 0.00947f
C49 a_18_1972# a_n33_639# 1.15e-19
C50 a_n76_4444# a_n33_3111# 1.15e-19
C51 a_n76_n4208# a_n33_n5541# 1.15e-19
C52 a_18_n5444# a_18_n6680# 0.00947f
C53 a_18_3208# w_n112_4344# 0.00199f
C54 w_n112_n5544# a_18_n4208# 0.00199f
C55 a_18_4444# a_n33_5583# 1.15e-19
C56 a_n33_6819# a_n33_8055# 0.0665f
C57 a_n33_n8013# a_n33_n9249# 0.0665f
C58 a_n33_n3069# a_18_n2972# 0.0417f
C59 a_n76_736# w_n112_n600# 0.00199f
C60 w_n112_n6780# a_n76_n7916# 0.00199f
C61 a_n33_n3069# w_n112_n1836# 4.13e-19
C62 w_n112_n8016# a_n33_n9249# 4.13e-19
C63 a_n33_n597# w_n112_n1836# 4.13e-19
C64 a_n76_6916# w_n112_8052# 0.00199f
C65 a_n76_n5444# a_n76_n4208# 0.00947f
C66 a_18_n5444# a_n33_n4305# 1.15e-19
C67 a_18_4444# a_n33_3111# 1.15e-19
C68 a_n33_n1833# a_n76_n1736# 0.0417f
C69 a_n33_n6777# a_18_n6680# 0.0417f
C70 a_18_736# a_18_n500# 0.00947f
C71 a_n33_n597# a_n76_n500# 0.0417f
C72 a_n76_n7916# a_n76_n9152# 0.00947f
C73 a_n33_n8013# a_18_n9152# 1.15e-19
C74 a_18_n7916# a_n33_n9249# 1.15e-19
C75 w_n112_n5544# a_n33_n5541# 0.106f
C76 a_18_n2972# w_n112_n1836# 0.00199f
C77 a_n76_n2972# w_n112_n3072# 0.0182f
C78 w_n112_n4308# a_n76_n2972# 0.00199f
C79 a_n76_6916# a_n33_8055# 1.15e-19
C80 a_n33_6819# a_n76_8152# 1.15e-19
C81 a_n33_n3069# a_n33_n4305# 0.0665f
C82 w_n112_n8016# a_18_n9152# 0.00199f
C83 w_n112_n9252# a_n76_n9152# 0.0182f
C84 a_18_n5444# a_18_n4208# 0.00947f
C85 a_n76_n500# w_n112_n1836# 0.00199f
C86 a_18_6916# w_n112_8052# 0.00199f
C87 a_n76_5680# w_n112_5580# 0.0182f
C88 a_n76_n1736# a_18_n1736# 0.747f
C89 w_n112_3108# a_n33_4347# 4.13e-19
C90 a_n33_3111# a_n76_3208# 0.0417f
C91 a_18_4444# a_18_3208# 0.00947f
C92 a_18_n7916# a_18_n9152# 0.00947f
C93 a_n33_639# a_n76_736# 0.0417f
C94 a_n76_5680# w_n112_6816# 0.00199f
C95 a_18_736# a_n33_1875# 1.15e-19
C96 a_n33_n6777# a_n33_n8013# 0.0665f
C97 w_n112_n5544# a_n76_n5444# 0.0182f
C98 a_n33_n597# a_18_n500# 0.0417f
C99 a_18_n2972# a_n33_n4305# 1.15e-19
C100 a_n33_n3069# a_18_n4208# 1.15e-19
C101 a_n76_n2972# a_n76_n4208# 0.00947f
C102 a_n76_6916# a_n76_8152# 0.00947f
C103 a_18_6916# a_n33_8055# 1.15e-19
C104 a_18_8152# w_n112_8052# 0.0182f
C105 w_n112_n8016# a_n33_n6777# 4.13e-19
C106 a_n76_n1736# w_n112_n600# 0.00199f
C107 a_18_n5444# a_n33_n5541# 0.0417f
C108 w_n112_636# a_18_736# 0.0182f
C109 w_n112_1872# a_18_736# 0.00199f
C110 a_18_n500# w_n112_n1836# 0.00199f
C111 a_n33_n9249# a_n76_n9152# 0.0417f
C112 a_18_5680# w_n112_5580# 0.0182f
C113 w_n112_3108# a_n76_4444# 0.00199f
C114 a_18_n6680# a_n33_n8013# 1.15e-19
C115 a_n33_n6777# a_18_n7916# 1.15e-19
C116 a_n76_n6680# a_n76_n7916# 0.00947f
C117 a_n76_3208# a_18_3208# 0.747f
C118 w_n112_n6780# a_18_n5444# 0.00199f
C119 a_n33_3111# a_18_3208# 0.0417f
C120 a_n33_n1833# a_n33_n3069# 0.0665f
C121 a_18_5680# w_n112_6816# 0.00199f
C122 a_18_8152# a_n33_8055# 0.0417f
C123 a_18_n2972# a_18_n4208# 0.00947f
C124 a_n76_n4208# w_n112_n3072# 0.00199f
C125 a_n33_6819# w_n112_5580# 4.13e-19
C126 a_n33_n597# a_n33_n1833# 0.0665f
C127 a_n76_n500# a_18_n500# 0.747f
C128 w_n112_n4308# a_n76_n4208# 0.0182f
C129 w_n112_n8016# a_18_n6680# 0.00199f
C130 a_n33_6819# w_n112_6816# 0.106f
C131 a_n76_n5444# a_18_n5444# 0.747f
C132 a_n76_n9152# a_18_n9152# 0.747f
C133 a_n33_n6777# a_n33_n5541# 0.0665f
C134 w_n112_636# a_n33_n597# 4.13e-19
C135 a_18_n6680# a_18_n7916# 0.00947f
C136 a_18_736# w_n112_n600# 0.00199f
C137 a_n33_n1833# a_18_n2972# 1.15e-19
C138 a_18_n1736# a_n33_n3069# 1.15e-19
C139 a_n76_n1736# a_n76_n2972# 0.00947f
C140 a_n33_n1833# w_n112_n1836# 0.106f
C141 a_n33_4347# w_n112_5580# 4.13e-19
C142 w_n112_3108# a_18_4444# 0.00199f
C143 w_n112_n6780# a_n33_n6777# 0.106f
C144 a_n76_3208# a_n33_1875# 1.15e-19
C145 w_n112_n5544# a_n76_n6680# 0.00199f
C146 a_n33_n597# a_18_n1736# 1.15e-19
C147 a_n76_5680# a_18_5680# 0.747f
C148 a_n33_3111# a_n33_1875# 0.0665f
C149 a_18_8152# a_n76_8152# 0.747f
C150 a_18_736# a_18_1972# 0.00947f
C151 a_n33_n4305# a_18_n4208# 0.0417f
C152 a_n76_n500# a_n33_n1833# 1.15e-19
C153 a_n76_6916# w_n112_5580# 0.00199f
C154 a_n76_5680# a_n33_6819# 1.15e-19
C155 w_n112_n8016# a_n33_n8013# 0.106f
C156 a_n76_6916# w_n112_6816# 0.0182f
C157 a_18_n6680# a_n33_n5541# 1.15e-19
C158 a_n76_n5444# a_n33_n6777# 1.15e-19
C159 a_18_n1736# a_18_n2972# 0.00947f
C160 a_18_n1736# w_n112_n1836# 0.0182f
C161 a_n76_n1736# w_n112_n3072# 0.00199f
C162 w_n112_636# a_n76_n500# 0.00199f
C163 a_n33_n597# w_n112_n600# 0.106f
C164 w_n112_1872# a_n76_3208# 0.00199f
C165 a_n33_n8013# a_18_n7916# 0.0417f
C166 w_n112_n6780# a_18_n6680# 0.0182f
C167 w_n112_1872# a_n33_3111# 4.13e-19
C168 w_n112_3108# a_n76_3208# 0.0182f
C169 a_n76_4444# w_n112_5580# 0.00199f
C170 w_n112_3108# a_n33_3111# 0.106f
C171 a_18_3208# a_n33_1875# 1.15e-19
C172 a_n76_3208# a_n76_1972# 0.00947f
C173 a_n76_5680# a_n33_4347# 1.15e-19
C174 a_n33_3111# a_n76_1972# 1.15e-19
C175 w_n112_n9252# a_n76_n7916# 0.00199f
C176 w_n112_n8016# a_18_n7916# 0.0182f
C177 a_18_736# a_n33_639# 0.0417f
C178 a_n33_n4305# a_n33_n5541# 0.0665f
C179 a_18_6916# w_n112_5580# 0.00199f
C180 a_18_n500# a_n33_n1833# 1.15e-19
C181 a_n76_5680# w_n112_4344# 0.00199f
C182 a_18_5680# a_n33_6819# 1.15e-19
C183 a_n76_5680# a_n76_6916# 0.00947f
C184 a_18_6916# w_n112_6816# 0.0182f
C185 w_n112_n5544# a_n76_n4208# 0.00199f
C186 a_n33_8055# w_n112_8052# 0.106f
C187 w_n112_636# a_18_n500# 0.00199f
C188 a_n33_n3069# a_n76_n2972# 0.0417f
C189 w_n112_1872# a_18_3208# 0.00199f
C190 a_n76_n500# w_n112_n600# 0.0182f
C191 w_n112_n6780# a_n33_n8013# 4.13e-19
C192 w_n112_n4308# a_18_n5444# 0.00199f
C193 w_n112_3108# a_18_3208# 0.0182f
C194 a_18_4444# w_n112_5580# 0.00199f
C195 a_18_n4208# a_n33_n5541# 1.15e-19
C196 a_n76_n5444# a_n33_n4305# 1.15e-19
C197 a_n76_5680# a_n76_4444# 0.00947f
C198 a_18_n500# a_18_n1736# 0.00947f
C199 a_18_5680# a_n33_4347# 1.15e-19
C200 a_18_8152# w_n112_6816# 0.00199f
C201 a_n33_3111# a_18_1972# 1.15e-19
C202 a_n33_n597# a_n33_639# 0.0665f
C203 a_18_736# a_n76_736# 0.747f
C204 a_n33_5583# w_n112_5580# 0.106f
C205 a_n33_n6777# a_n76_n6680# 0.0417f
C206 a_18_5680# w_n112_4344# 0.00199f
C207 a_n76_n7916# a_n33_n9249# 1.15e-19
C208 a_n33_n8013# a_n76_n9152# 1.15e-19
C209 a_n33_5583# w_n112_6816# 4.13e-19
C210 a_n76_n2972# a_18_n2972# 0.747f
C211 a_n33_n3069# w_n112_n3072# 0.106f
C212 a_n76_n2972# w_n112_n1836# 0.00199f
C213 w_n112_n6780# a_18_n7916# 0.00199f
C214 w_n112_n4308# a_n33_n3069# 4.13e-19
C215 w_n112_636# a_n33_1875# 4.13e-19
C216 a_n76_8152# w_n112_8052# 0.0182f
C217 a_n33_6819# a_n76_6916# 0.0417f
C218 w_n112_n9252# a_n33_n9249# 0.106f
C219 w_n112_n8016# a_n76_n9152# 0.00199f
C220 a_18_n500# w_n112_n600# 0.0182f
C221 w_n112_1872# a_n33_1875# 0.106f
C222 w_n112_3108# a_n33_1875# 4.13e-19
C223 a_n33_1875# a_n76_1972# 0.0417f
C224 a_18_3208# a_18_1972# 0.00947f
C225 a_n33_n1833# a_18_n1736# 0.0417f
C226 a_n76_n6680# a_18_n6680# 0.747f
C227 a_n33_n597# a_n76_736# 1.15e-19
C228 a_n76_n500# a_n33_639# 1.15e-19
C229 a_n33_8055# a_n76_8152# 0.0417f
C230 w_n112_n6780# a_n33_n5541# 4.13e-19
C231 a_18_n2972# w_n112_n3072# 0.0182f
C232 w_n112_n4308# a_18_n2972# 0.00199f
C233 a_n33_4347# w_n112_4344# 0.106f
C234 a_18_5680# a_18_6916# 0.00947f
C235 a_n76_5680# a_n33_5583# 0.0417f
C236 a_n33_n3069# a_n76_n4208# 1.15e-19
C237 a_n76_n2972# a_n33_n4305# 1.15e-19
C238 w_n112_n9252# a_18_n9152# 0.0182f
C239 w_n112_636# a_n76_1972# 0.00199f
C240 a_n33_6819# a_18_6916# 0.0417f
C241 a_n33_n1833# w_n112_n600# 4.13e-19
C242 w_n112_1872# a_n76_1972# 0.0182f
C243 a_n76_n5444# a_n33_n5541# 0.0417f
C244 w_n112_3108# a_n76_1972# 0.00199f
C245 a_n33_1875# a_18_1972# 0.0417f
C246 a_18_5680# a_18_4444# 0.00947f
C247 a_n33_4347# a_n76_4444# 0.0417f
C248 a_n76_n6680# a_n33_n8013# 1.15e-19
C249 a_n33_n6777# a_n76_n7916# 1.15e-19
C250 w_n112_n5544# a_18_n5444# 0.0182f
C251 w_n112_n6780# a_n76_n5444# 0.00199f
C252 a_18_n500# a_n33_639# 1.15e-19
C253 a_n76_n500# a_n76_736# 0.00947f
C254 a_18_8152# a_n33_6819# 1.15e-19
C255 a_n33_n4305# w_n112_n3072# 4.13e-19
C256 a_n76_4444# w_n112_4344# 0.0182f
C257 w_n112_n4308# a_n33_n4305# 0.106f
C258 a_18_5680# a_n33_5583# 0.0417f
C259 w_n112_n8016# a_n76_n6680# 0.00199f
C260 a_18_n1736# w_n112_n600# 0.00199f
C261 w_n112_636# a_18_1972# 0.00199f
C262 a_n33_6819# a_n33_5583# 0.0665f
C263 a_n76_6916# a_18_6916# 0.747f
C264 w_n112_1872# a_18_1972# 0.0182f
C265 a_n33_n9249# a_18_n9152# 0.0417f
C266 w_n112_3108# a_18_1972# 0.00199f
C267 a_n33_n1833# a_n76_n2972# 1.15e-19
C268 a_n76_n1736# a_n33_n3069# 1.15e-19
C269 a_n76_1972# a_18_1972# 0.747f
C270 a_n33_1875# a_n33_639# 0.0665f
C271 a_n33_4347# a_18_4444# 0.0417f
C272 a_18_n9152# VSUBS 0.426f
C273 a_n76_n9152# VSUBS 0.426f
C274 a_n33_n9249# VSUBS 0.192f
C275 a_18_n7916# VSUBS 0.415f
C276 a_n76_n7916# VSUBS 0.415f
C277 a_n33_n8013# VSUBS 0.156f
C278 a_18_n6680# VSUBS 0.415f
C279 a_n76_n6680# VSUBS 0.415f
C280 a_n33_n6777# VSUBS 0.156f
C281 a_18_n5444# VSUBS 0.415f
C282 a_n76_n5444# VSUBS 0.415f
C283 a_n33_n5541# VSUBS 0.156f
C284 a_18_n4208# VSUBS 0.415f
C285 a_n76_n4208# VSUBS 0.415f
C286 a_n33_n4305# VSUBS 0.156f
C287 a_18_n2972# VSUBS 0.415f
C288 a_n76_n2972# VSUBS 0.415f
C289 a_n33_n3069# VSUBS 0.156f
C290 a_18_n1736# VSUBS 0.415f
C291 a_n76_n1736# VSUBS 0.415f
C292 a_n33_n1833# VSUBS 0.156f
C293 a_18_n500# VSUBS 0.415f
C294 a_n76_n500# VSUBS 0.415f
C295 a_n33_n597# VSUBS 0.156f
C296 a_18_736# VSUBS 0.415f
C297 a_n76_736# VSUBS 0.415f
C298 a_n33_639# VSUBS 0.156f
C299 a_18_1972# VSUBS 0.415f
C300 a_n76_1972# VSUBS 0.415f
C301 a_n33_1875# VSUBS 0.156f
C302 a_18_3208# VSUBS 0.415f
C303 a_n76_3208# VSUBS 0.415f
C304 a_n33_3111# VSUBS 0.156f
C305 a_18_4444# VSUBS 0.415f
C306 a_n76_4444# VSUBS 0.415f
C307 a_n33_4347# VSUBS 0.156f
C308 a_18_5680# VSUBS 0.415f
C309 a_n76_5680# VSUBS 0.415f
C310 a_n33_5583# VSUBS 0.156f
C311 a_18_6916# VSUBS 0.415f
C312 a_n76_6916# VSUBS 0.415f
C313 a_n33_6819# VSUBS 0.156f
C314 a_18_8152# VSUBS 0.426f
C315 a_n76_8152# VSUBS 0.426f
C316 a_n33_8055# VSUBS 0.192f
C317 w_n112_n9252# VSUBS 0.806f
C318 w_n112_n8016# VSUBS 0.806f
C319 w_n112_n6780# VSUBS 0.806f
C320 w_n112_n5544# VSUBS 0.806f
C321 w_n112_n4308# VSUBS 0.806f
C322 w_n112_n3072# VSUBS 0.806f
C323 w_n112_n1836# VSUBS 0.806f
C324 w_n112_n600# VSUBS 0.806f
C325 w_n112_636# VSUBS 0.806f
C326 w_n112_1872# VSUBS 0.806f
C327 w_n112_3108# VSUBS 0.806f
C328 w_n112_4344# VSUBS 0.806f
C329 w_n112_5580# VSUBS 0.806f
C330 w_n112_6816# VSUBS 0.806f
C331 w_n112_8052# VSUBS 0.806f
.ends

.subckt sky130_fd_pr__nfet_01v8_MHE452 a_n158_n359# a_n100_957# a_100_n1295# a_n158_577#
+ a_n100_21# a_100_109# a_n100_n915# a_100_n827# a_n100_489# a_100_1045# a_n158_n1295#
+ a_n158_n827# a_100_577# a_n158_1045# a_n100_n447# a_n158_109# a_100_n359# a_n100_n1383#
+ VSUBS
X0 a_100_n827# a_n100_n915# a_n158_n827# VSUBS sky130_fd_pr__nfet_01v8 ad=0.363 pd=3.08 as=0.363 ps=3.08 w=1.25 l=1
**devattr s=14500,616 d=14500,616
X1 a_100_n359# a_n100_n447# a_n158_n359# VSUBS sky130_fd_pr__nfet_01v8 ad=0.363 pd=3.08 as=0.363 ps=3.08 w=1.25 l=1
**devattr s=14500,616 d=14500,616
X2 a_100_577# a_n100_489# a_n158_577# VSUBS sky130_fd_pr__nfet_01v8 ad=0.363 pd=3.08 as=0.363 ps=3.08 w=1.25 l=1
**devattr s=14500,616 d=14500,616
X3 a_100_1045# a_n100_957# a_n158_1045# VSUBS sky130_fd_pr__nfet_01v8 ad=0.363 pd=3.08 as=0.363 ps=3.08 w=1.25 l=1
**devattr s=14500,616 d=14500,616
X4 a_100_n1295# a_n100_n1383# a_n158_n1295# VSUBS sky130_fd_pr__nfet_01v8 ad=0.363 pd=3.08 as=0.363 ps=3.08 w=1.25 l=1
**devattr s=14500,616 d=14500,616
X5 a_100_109# a_n100_21# a_n158_109# VSUBS sky130_fd_pr__nfet_01v8 ad=0.363 pd=3.08 as=0.363 ps=3.08 w=1.25 l=1
**devattr s=14500,616 d=14500,616
C0 a_100_n359# a_n100_n447# 0.0322f
C1 a_n100_957# a_n158_1045# 0.0322f
C2 a_n158_n827# a_100_n827# 0.0693f
C3 a_n158_n359# a_n158_n827# 0.0113f
C4 a_n100_n1383# a_n100_n915# 0.205f
C5 a_n158_1045# a_100_1045# 0.0693f
C6 a_n158_n827# a_n100_n915# 0.0322f
C7 a_n100_957# a_n100_489# 0.205f
C8 a_100_n359# a_100_109# 0.0113f
C9 a_n100_n915# a_100_n827# 0.0322f
C10 a_n158_1045# a_n158_577# 0.0113f
C11 a_100_n1295# a_n158_n1295# 0.0693f
C12 a_100_1045# a_100_577# 0.0113f
C13 a_n158_n359# a_n100_n447# 0.0322f
C14 a_n158_n359# a_n158_109# 0.0113f
C15 a_n100_21# a_n100_489# 0.205f
C16 a_n100_489# a_n158_577# 0.0322f
C17 a_n100_n1383# a_100_n1295# 0.0322f
C18 a_n100_n447# a_n100_n915# 0.205f
C19 a_n158_577# a_100_577# 0.0693f
C20 a_100_577# a_100_109# 0.0113f
C21 a_100_n1295# a_100_n827# 0.0113f
C22 a_n100_957# a_100_1045# 0.0322f
C23 a_n100_n447# a_n100_21# 0.205f
C24 a_n100_n1383# a_n158_n1295# 0.0322f
C25 a_n158_109# a_n100_21# 0.0322f
C26 a_100_n359# a_100_n827# 0.0113f
C27 a_n158_109# a_n158_577# 0.0113f
C28 a_100_n359# a_n158_n359# 0.0693f
C29 a_n158_109# a_100_109# 0.0693f
C30 a_n158_n827# a_n158_n1295# 0.0113f
C31 a_n100_489# a_100_577# 0.0322f
C32 a_n100_21# a_100_109# 0.0322f
C33 a_100_n1295# VSUBS 0.14f
C34 a_n158_n1295# VSUBS 0.14f
C35 a_n100_n1383# VSUBS 0.553f
C36 a_100_n827# VSUBS 0.13f
C37 a_n158_n827# VSUBS 0.13f
C38 a_n100_n915# VSUBS 0.441f
C39 a_100_n359# VSUBS 0.13f
C40 a_n158_n359# VSUBS 0.13f
C41 a_n100_n447# VSUBS 0.441f
C42 a_100_109# VSUBS 0.13f
C43 a_n158_109# VSUBS 0.13f
C44 a_n100_21# VSUBS 0.441f
C45 a_100_577# VSUBS 0.13f
C46 a_n158_577# VSUBS 0.13f
C47 a_n100_489# VSUBS 0.441f
C48 a_100_1045# VSUBS 0.14f
C49 a_n158_1045# VSUBS 0.14f
C50 a_n100_957# VSUBS 0.553f
.ends

.subckt sky130_fd_pr__pfet_01v8_P2UXFR a_n300_n1215# w_n394_n1218# a_n358_n1118# a_n300_21#
+ a_300_118# w_n394_18# a_300_n1118# a_n358_118# VSUBS
X0 a_300_118# a_n300_21# a_n358_118# w_n394_18# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=3
**devattr s=58000,2116 d=58000,2116
X1 a_300_n1118# a_n300_n1215# a_n358_n1118# w_n394_n1218# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=3
**devattr s=58000,2116 d=58000,2116
C0 w_n394_18# a_300_118# 0.0187f
C1 a_n358_n1118# a_300_n1118# 0.107f
C2 a_n358_118# a_n300_21# 0.184f
C3 a_n358_n1118# a_n358_118# 0.0105f
C4 w_n394_n1218# a_n300_21# 0.00346f
C5 a_n358_n1118# w_n394_n1218# 0.0187f
C6 w_n394_18# a_300_n1118# 0.0023f
C7 a_n358_118# w_n394_18# 0.0187f
C8 w_n394_18# a_n300_21# 0.382f
C9 a_n358_n1118# w_n394_18# 0.0023f
C10 a_n300_n1215# a_300_n1118# 0.184f
C11 w_n394_n1218# a_n300_n1215# 0.382f
C12 a_n300_n1215# a_n300_21# 0.62f
C13 a_n358_n1118# a_n300_n1215# 0.184f
C14 w_n394_18# a_n300_n1215# 0.00346f
C15 a_300_n1118# a_300_118# 0.0105f
C16 a_n358_118# a_300_118# 0.107f
C17 w_n394_n1218# a_300_118# 0.0023f
C18 a_n300_21# a_300_118# 0.184f
C19 w_n394_n1218# a_300_n1118# 0.0187f
C20 a_n358_118# w_n394_n1218# 0.0023f
C21 a_300_n1118# VSUBS 0.536f
C22 a_n358_n1118# VSUBS 0.536f
C23 a_n300_n1215# VSUBS 1.08f
C24 a_300_118# VSUBS 0.536f
C25 a_n358_118# VSUBS 0.536f
C26 a_n300_21# VSUBS 1.08f
C27 w_n394_n1218# VSUBS 2.84f
C28 w_n394_18# VSUBS 2.84f
.ends

.subckt sky130_fd_pr__pfet_01v8_MGA63L a_18_n500# a_n33_n597# w_n112_n600# a_n76_n500#
+ VSUBS
X0 a_18_n500# a_n33_n597# a_n76_n500# w_n112_n600# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
C0 w_n112_n600# a_n33_n597# 0.106f
C1 a_18_n500# a_n33_n597# 0.0417f
C2 w_n112_n600# a_18_n500# 0.0182f
C3 a_n76_n500# a_n33_n597# 0.0417f
C4 w_n112_n600# a_n76_n500# 0.0182f
C5 a_18_n500# a_n76_n500# 0.747f
C6 a_18_n500# VSUBS 0.437f
C7 a_n76_n500# VSUBS 0.437f
C8 a_n33_n597# VSUBS 0.228f
C9 w_n112_n600# VSUBS 0.806f
.ends

.subckt sky130_fd_pr__nfet_01v8_VT3ZQW a_n158_n125# a_n100_n213# a_100_n125# VSUBS
X0 a_100_n125# a_n100_n213# a_n158_n125# VSUBS sky130_fd_pr__nfet_01v8 ad=0.363 pd=3.08 as=0.363 ps=3.08 w=1.25 l=1
**devattr s=14500,616 d=14500,616
C0 a_n100_n213# a_n158_n125# 0.0322f
C1 a_100_n125# a_n158_n125# 0.0693f
C2 a_n100_n213# a_100_n125# 0.0322f
C3 a_100_n125# VSUBS 0.151f
C4 a_n158_n125# VSUBS 0.151f
C5 a_n100_n213# VSUBS 0.664f
.ends

.subckt sky130_fd_pr__pfet_01v8_RRUZAE a_n358_n2972# a_n300_n1833# a_n300_n3069# w_n394_n1836#
+ w_n394_1872# a_n358_n1736# a_300_736# a_300_1972# a_300_n2972# w_n394_636# w_n394_n3072#
+ a_n300_n597# a_300_n500# a_n300_639# a_n358_1972# a_n300_1875# w_n394_n600# a_300_n1736#
+ a_n358_n500# a_n358_736# VSUBS
X0 a_300_n500# a_n300_n597# a_n358_n500# w_n394_n600# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=3
**devattr s=58000,2116 d=58000,2116
X1 a_300_736# a_n300_639# a_n358_736# w_n394_636# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=3
**devattr s=58000,2116 d=58000,2116
X2 a_300_n2972# a_n300_n3069# a_n358_n2972# w_n394_n3072# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=3
**devattr s=58000,2116 d=58000,2116
X3 a_300_1972# a_n300_1875# a_n358_1972# w_n394_1872# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=3
**devattr s=58000,2116 d=58000,2116
X4 a_300_n1736# a_n300_n1833# a_n358_n1736# w_n394_n1836# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=3
**devattr s=58000,2116 d=58000,2116
C0 a_n358_736# a_n358_1972# 0.0105f
C1 a_n300_639# a_n300_n597# 0.62f
C2 a_n300_639# a_n300_1875# 0.62f
C3 a_300_1972# w_n394_636# 0.0023f
C4 a_300_n500# w_n394_636# 0.0023f
C5 a_n358_n500# a_300_n500# 0.107f
C6 a_300_736# a_300_1972# 0.0105f
C7 a_n300_n1833# a_n300_n597# 0.62f
C8 a_n358_n1736# a_300_n1736# 0.107f
C9 w_n394_1872# a_300_736# 0.0023f
C10 a_n358_n2972# w_n394_n1836# 0.0023f
C11 a_300_736# a_300_n500# 0.0105f
C12 w_n394_n1836# a_n300_n1833# 0.382f
C13 a_300_n2972# w_n394_n3072# 0.0187f
C14 a_n300_1875# a_n358_1972# 0.184f
C15 a_n358_736# w_n394_636# 0.0187f
C16 a_n358_n500# a_n358_736# 0.0105f
C17 w_n394_1872# a_300_1972# 0.0187f
C18 a_300_736# a_n358_736# 0.107f
C19 a_n300_639# w_n394_n600# 0.00346f
C20 w_n394_n1836# a_n300_n3069# 0.00346f
C21 a_n358_n1736# w_n394_n1836# 0.0187f
C22 a_n300_n597# w_n394_636# 0.00346f
C23 a_n358_n500# a_n300_n597# 0.184f
C24 a_n300_1875# w_n394_636# 0.00346f
C25 w_n394_1872# a_n358_736# 0.0023f
C26 w_n394_n600# a_n300_n1833# 0.00346f
C27 a_n358_n500# w_n394_n1836# 0.0023f
C28 a_300_n500# a_300_n1736# 0.0105f
C29 a_n358_n2972# w_n394_n3072# 0.0187f
C30 a_n300_n1833# w_n394_n3072# 0.00346f
C31 a_n300_1875# a_300_1972# 0.184f
C32 a_n358_n1736# w_n394_n600# 0.0023f
C33 a_n300_n597# a_300_n500# 0.184f
C34 w_n394_1872# a_n300_1875# 0.382f
C35 a_n300_n3069# w_n394_n3072# 0.382f
C36 a_n358_n2972# a_300_n2972# 0.107f
C37 a_n358_n1736# w_n394_n3072# 0.0023f
C38 w_n394_n1836# a_300_n500# 0.0023f
C39 a_n358_n500# w_n394_n600# 0.0187f
C40 a_300_736# w_n394_n600# 0.0023f
C41 w_n394_n1836# a_300_n1736# 0.0187f
C42 a_300_n2972# a_n300_n3069# 0.184f
C43 w_n394_n600# a_300_n500# 0.0187f
C44 w_n394_n1836# a_n300_n597# 0.00346f
C45 a_n358_736# w_n394_n600# 0.0023f
C46 w_n394_n600# a_300_n1736# 0.0023f
C47 a_n358_n2972# a_n300_n3069# 0.184f
C48 a_n300_639# w_n394_636# 0.382f
C49 a_n358_n2972# a_n358_n1736# 0.0105f
C50 a_n300_n1833# a_n300_n3069# 0.62f
C51 a_300_n1736# w_n394_n3072# 0.0023f
C52 a_n358_n1736# a_n300_n1833# 0.184f
C53 a_n300_639# a_300_736# 0.184f
C54 w_n394_n600# a_n300_n597# 0.382f
C55 w_n394_636# a_n358_1972# 0.0023f
C56 a_300_n2972# a_300_n1736# 0.0105f
C57 a_n300_639# w_n394_1872# 0.00346f
C58 a_n358_n500# a_n358_n1736# 0.0105f
C59 a_n300_639# a_n358_736# 0.184f
C60 a_300_1972# a_n358_1972# 0.107f
C61 a_n358_n500# w_n394_636# 0.0023f
C62 w_n394_1872# a_n358_1972# 0.0187f
C63 a_300_n2972# w_n394_n1836# 0.0023f
C64 a_300_736# w_n394_636# 0.0187f
C65 a_n300_n1833# a_300_n1736# 0.184f
C66 a_300_n2972# VSUBS 0.536f
C67 a_n358_n2972# VSUBS 0.536f
C68 a_n300_n3069# VSUBS 1.08f
C69 a_300_n1736# VSUBS 0.524f
C70 a_n358_n1736# VSUBS 0.524f
C71 a_n300_n1833# VSUBS 0.739f
C72 a_300_n500# VSUBS 0.524f
C73 a_n358_n500# VSUBS 0.524f
C74 a_n300_n597# VSUBS 0.739f
C75 a_300_736# VSUBS 0.524f
C76 a_n358_736# VSUBS 0.524f
C77 a_n300_639# VSUBS 0.739f
C78 a_300_1972# VSUBS 0.536f
C79 a_n358_1972# VSUBS 0.536f
C80 a_n300_1875# VSUBS 1.08f
C81 w_n394_n3072# VSUBS 2.84f
C82 w_n394_n1836# VSUBS 2.84f
C83 w_n394_n600# VSUBS 2.84f
C84 w_n394_636# VSUBS 2.84f
C85 w_n394_1872# VSUBS 2.84f
.ends

.subckt sky130_fd_pr__pfet_01v8_8DHNHY w_n112_636# a_n33_n5541# a_n33_n8013# a_n76_736#
+ a_n33_9291# w_n112_1872# a_18_9388# w_n112_4344# a_18_n500# a_18_n2972# a_18_n5444#
+ a_n76_n1736# a_n33_3111# a_n76_n4208# a_18_3208# w_n112_9288# a_n76_n7916# a_n33_n1833#
+ a_18_6916# a_n76_5680# w_n112_n3072# a_n76_n10388# a_n33_n4305# a_n33_5583# a_n76_8152#
+ w_n112_n6780# a_n33_8055# a_n33_n3069# a_n33_639# w_n112_n9252# w_n112_3108# a_18_n10388#
+ w_n112_6816# a_n33_n6777# a_n33_n597# w_n112_n10488# a_n33_n9249# a_18_n1736# a_18_n4208#
+ a_18_n7916# a_n76_1972# a_n33_1875# w_n112_n600# a_n76_n6680# a_18_736# a_n76_4444#
+ a_18_5680# a_n33_4347# w_n112_n5544# a_n76_n9152# a_18_8152# w_n112_n8016# a_n76_n500#
+ a_n76_9388# w_n112_5580# w_n112_8052# a_18_n6680# a_n76_n2972# a_18_1972# a_n76_3208#
+ a_n76_n5444# a_18_4444# a_n76_6916# w_n112_n1836# a_n33_n10485# a_18_n9152# a_n33_6819#
+ w_n112_n4308# VSUBS
X0 a_18_3208# a_n33_3111# a_n76_3208# w_n112_3108# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X1 a_18_n6680# a_n33_n6777# a_n76_n6680# w_n112_n6780# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X2 a_18_9388# a_n33_9291# a_n76_9388# w_n112_9288# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X3 a_18_n500# a_n33_n597# a_n76_n500# w_n112_n600# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X4 a_18_n9152# a_n33_n9249# a_n76_n9152# w_n112_n9252# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X5 a_18_736# a_n33_639# a_n76_736# w_n112_636# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X6 a_18_n2972# a_n33_n3069# a_n76_n2972# w_n112_n3072# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X7 a_18_n7916# a_n33_n8013# a_n76_n7916# w_n112_n8016# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X8 a_18_5680# a_n33_5583# a_n76_5680# w_n112_5580# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X9 a_18_n5444# a_n33_n5541# a_n76_n5444# w_n112_n5544# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X10 a_18_8152# a_n33_8055# a_n76_8152# w_n112_8052# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X11 a_18_n1736# a_n33_n1833# a_n76_n1736# w_n112_n1836# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X12 a_18_6916# a_n33_6819# a_n76_6916# w_n112_6816# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X13 a_18_1972# a_n33_1875# a_n76_1972# w_n112_1872# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X14 a_18_n4208# a_n33_n4305# a_n76_n4208# w_n112_n4308# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X15 a_18_4444# a_n33_4347# a_n76_4444# w_n112_4344# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
X16 a_18_n10388# a_n33_n10485# a_n76_n10388# w_n112_n10488# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=0.18
**devattr s=58000,2116 d=58000,2116
C0 a_n33_4347# a_n33_3111# 0.0665f
C1 w_n112_4344# a_n33_5583# 4.13e-19
C2 a_n33_n8013# w_n112_n9252# 4.13e-19
C3 a_n76_n6680# a_n76_n7916# 0.00947f
C4 a_18_n6680# a_n33_n8013# 1.15e-19
C5 w_n112_n8016# a_n76_n9152# 0.00199f
C6 a_n33_9291# a_n76_8152# 1.15e-19
C7 a_18_n500# w_n112_n600# 0.0182f
C8 a_n76_n500# a_n33_n1833# 1.15e-19
C9 a_18_n9152# w_n112_n9252# 0.0182f
C10 a_n76_n1736# a_18_n1736# 0.747f
C11 a_n33_4347# w_n112_5580# 4.13e-19
C12 a_n76_5680# w_n112_5580# 0.0182f
C13 a_n33_9291# a_n76_9388# 0.0417f
C14 a_n33_n3069# a_18_n2972# 0.0417f
C15 w_n112_1872# a_n33_639# 4.13e-19
C16 a_n33_n9249# a_n33_n8013# 0.0665f
C17 w_n112_n6780# a_n33_n8013# 4.13e-19
C18 a_18_3208# w_n112_3108# 0.0182f
C19 a_n76_n5444# a_18_n5444# 0.747f
C20 w_n112_n8016# a_n76_n7916# 0.0182f
C21 w_n112_n5544# a_n33_n6777# 4.13e-19
C22 a_n33_n9249# a_18_n9152# 0.0417f
C23 a_n33_n9249# w_n112_n10488# 4.13e-19
C24 w_n112_636# a_n33_639# 0.106f
C25 a_n33_n597# a_n33_639# 0.0665f
C26 a_18_n4208# a_n76_n4208# 0.747f
C27 a_n33_n1833# w_n112_n600# 4.13e-19
C28 a_18_n500# a_n33_n1833# 1.15e-19
C29 a_n33_1875# a_n76_1972# 0.0417f
C30 a_18_3208# a_18_1972# 0.00947f
C31 a_n33_5583# w_n112_5580# 0.106f
C32 a_n33_n10485# w_n112_n9252# 4.13e-19
C33 a_n76_8152# w_n112_6816# 0.00199f
C34 a_n33_n1833# a_n76_n2972# 1.15e-19
C35 a_18_9388# w_n112_9288# 0.0182f
C36 a_n76_n1736# a_n33_n3069# 1.15e-19
C37 a_n76_n9152# a_n76_n7916# 0.00947f
C38 a_18_n9152# a_n33_n8013# 1.15e-19
C39 a_n33_n3069# a_n33_n4305# 0.0665f
C40 a_n76_3208# a_18_3208# 0.747f
C41 w_n112_n4308# a_18_n4208# 0.0182f
C42 w_n112_n5544# a_18_n6680# 0.00199f
C43 w_n112_1872# a_n33_3111# 4.13e-19
C44 w_n112_1872# a_n76_736# 0.00199f
C45 a_18_n4208# a_n33_n5541# 1.15e-19
C46 a_18_n9152# w_n112_n10488# 0.00199f
C47 a_n33_1875# w_n112_3108# 4.13e-19
C48 a_n33_n5541# a_n76_n6680# 1.15e-19
C49 a_n76_n5444# a_n33_n6777# 1.15e-19
C50 a_18_6916# w_n112_6816# 0.0182f
C51 a_n33_n9249# a_n33_n10485# 0.0665f
C52 w_n112_n8016# a_18_n7916# 0.0182f
C53 w_n112_636# a_n76_736# 0.0182f
C54 a_n76_5680# a_n33_6819# 1.15e-19
C55 a_n76_n500# a_n33_639# 1.15e-19
C56 a_n33_n597# a_n76_736# 1.15e-19
C57 a_18_n10388# w_n112_n9252# 0.00199f
C58 w_n112_9288# a_18_8152# 0.00199f
C59 a_18_6916# a_n33_5583# 1.15e-19
C60 w_n112_3108# a_n76_1972# 0.00199f
C61 w_n112_n1836# a_18_n1736# 0.0182f
C62 a_n33_1875# a_18_1972# 0.0417f
C63 a_n76_n2972# a_n76_n4208# 0.00947f
C64 a_18_n2972# a_n33_n4305# 1.15e-19
C65 a_n33_6819# w_n112_6816# 0.106f
C66 a_18_n4208# a_18_n5444# 0.00947f
C67 a_n33_8055# w_n112_9288# 4.13e-19
C68 a_18_4444# a_n33_4347# 0.0417f
C69 a_n33_n597# a_18_n1736# 1.15e-19
C70 a_18_3208# w_n112_4344# 0.00199f
C71 a_n76_3208# a_n33_1875# 1.15e-19
C72 w_n112_8052# a_18_9388# 0.00199f
C73 a_n76_n9152# a_n76_n10388# 0.00947f
C74 a_18_n9152# a_n33_n10485# 1.15e-19
C75 a_n33_n9249# a_18_n10388# 1.15e-19
C76 w_n112_1872# a_18_736# 0.00199f
C77 a_18_n4208# w_n112_n3072# 0.00199f
C78 a_n33_n10485# w_n112_n10488# 0.106f
C79 w_n112_n4308# a_n76_n2972# 0.00199f
C80 a_n76_1972# a_18_1972# 0.747f
C81 a_n33_5583# a_n33_6819# 0.0665f
C82 w_n112_636# a_18_736# 0.0182f
C83 w_n112_n600# a_n33_639# 4.13e-19
C84 a_n76_n500# a_n76_736# 0.00947f
C85 a_n33_n597# a_18_736# 1.15e-19
C86 a_18_n500# a_n33_639# 1.15e-19
C87 a_n76_3208# a_n76_1972# 0.00947f
C88 w_n112_n6780# a_n76_n5444# 0.00199f
C89 a_18_n7916# a_n76_n7916# 0.747f
C90 a_n76_9388# a_18_9388# 0.747f
C91 a_18_4444# a_n33_5583# 1.15e-19
C92 w_n112_3108# a_18_1972# 0.00199f
C93 w_n112_n1836# a_n33_n3069# 4.13e-19
C94 w_n112_4344# a_18_5680# 0.00199f
C95 a_18_3208# a_n33_3111# 0.0417f
C96 a_n33_1875# a_n33_639# 0.0665f
C97 w_n112_8052# a_18_8152# 0.0182f
C98 a_18_n9152# a_18_n10388# 0.00947f
C99 a_n76_5680# a_n33_4347# 1.15e-19
C100 a_n76_3208# w_n112_3108# 0.0182f
C101 a_18_n10388# w_n112_n10488# 0.0182f
C102 w_n112_5580# a_n76_6916# 0.00199f
C103 a_n33_n6777# a_n76_n6680# 0.0417f
C104 w_n112_8052# a_n33_8055# 0.106f
C105 w_n112_8052# a_n76_6916# 0.00199f
C106 w_n112_n5544# a_n33_n4305# 4.13e-19
C107 a_18_8152# a_n76_8152# 0.747f
C108 a_n76_4444# w_n112_3108# 0.00199f
C109 a_n76_1972# a_n33_639# 1.15e-19
C110 a_n76_5680# w_n112_6816# 0.00199f
C111 a_n76_n2972# w_n112_n3072# 0.0182f
C112 a_n33_8055# a_n76_8152# 0.0417f
C113 a_n76_6916# a_n76_8152# 0.00947f
C114 w_n112_n1836# a_18_n2972# 0.00199f
C115 w_n112_n600# a_n76_736# 0.00199f
C116 a_18_6916# a_18_8152# 0.00947f
C117 w_n112_n8016# a_n33_n6777# 4.13e-19
C118 a_n76_9388# a_n33_8055# 1.15e-19
C119 a_n76_5680# a_n33_5583# 0.0417f
C120 a_n33_5583# a_n33_4347# 0.0665f
C121 a_n33_1875# a_n33_3111# 0.0665f
C122 a_n33_1875# a_n76_736# 1.15e-19
C123 a_18_6916# a_n33_8055# 1.15e-19
C124 a_n76_n6680# a_18_n6680# 0.747f
C125 a_n33_n10485# a_18_n10388# 0.0417f
C126 a_18_6916# a_n76_6916# 0.747f
C127 a_18_5680# w_n112_5580# 0.0182f
C128 a_18_n4208# a_n33_n3069# 1.15e-19
C129 a_18_n1736# w_n112_n600# 0.00199f
C130 a_18_n500# a_18_n1736# 0.00947f
C131 w_n112_n4308# a_n76_n4208# 0.0182f
C132 a_n33_5583# w_n112_6816# 4.13e-19
C133 a_n33_9291# a_18_9388# 0.0417f
C134 a_n76_3208# a_n76_4444# 0.00947f
C135 a_n33_n5541# a_n76_n4208# 1.15e-19
C136 a_n76_n5444# a_n33_n4305# 1.15e-19
C137 a_18_8152# a_n33_6819# 1.15e-19
C138 a_n33_n1833# w_n112_n3072# 4.13e-19
C139 a_n33_3111# a_n76_1972# 1.15e-19
C140 a_18_1972# a_n33_639# 1.15e-19
C141 a_n76_1972# a_n76_736# 0.00947f
C142 w_n112_n6780# a_n76_n6680# 0.0182f
C143 a_n76_n1736# w_n112_n1836# 0.0182f
C144 a_n33_8055# a_n33_6819# 0.0665f
C145 w_n112_n8016# a_18_n6680# 0.00199f
C146 w_n112_n5544# a_n76_n5444# 0.0182f
C147 a_n76_6916# a_n33_6819# 0.0417f
C148 w_n112_n600# a_18_736# 0.00199f
C149 a_18_n500# a_18_736# 0.00947f
C150 w_n112_n4308# a_n33_n5541# 4.13e-19
C151 a_n33_n597# a_n76_n1736# 1.15e-19
C152 w_n112_3108# a_n33_3111# 0.106f
C153 a_18_n4208# a_18_n2972# 0.00947f
C154 a_n76_3208# w_n112_4344# 0.00199f
C155 a_n33_1875# a_18_736# 1.15e-19
C156 a_18_6916# a_18_5680# 0.00947f
C157 a_n76_n6680# a_n33_n8013# 1.15e-19
C158 a_n33_n6777# a_n76_n7916# 1.15e-19
C159 w_n112_n8016# a_n33_n9249# 4.13e-19
C160 a_n33_9291# a_18_8152# 1.15e-19
C161 a_n76_n9152# w_n112_n9252# 0.0182f
C162 a_n33_n1833# a_18_n1736# 0.0417f
C163 w_n112_4344# a_n76_4444# 0.0182f
C164 a_n33_9291# a_n33_8055# 0.0665f
C165 a_18_3208# a_18_4444# 0.00947f
C166 a_n76_n4208# w_n112_n3072# 0.00199f
C167 a_n33_n3069# a_n76_n2972# 0.0417f
C168 a_n33_3111# a_18_1972# 1.15e-19
C169 w_n112_n4308# a_18_n5444# 0.00199f
C170 a_n33_n5541# a_18_n5444# 0.0417f
C171 a_18_5680# a_n33_6819# 1.15e-19
C172 w_n112_n8016# a_n33_n8013# 0.106f
C173 a_n33_n9249# a_n76_n9152# 0.0417f
C174 a_n76_n7916# w_n112_n9252# 0.00199f
C175 a_n76_3208# a_n33_3111# 0.0417f
C176 w_n112_n8016# a_18_n9152# 0.00199f
C177 a_n76_n500# a_n76_n1736# 0.00947f
C178 a_18_n4208# a_n33_n4305# 0.0417f
C179 a_n76_4444# a_n33_3111# 1.15e-19
C180 a_18_4444# a_18_5680# 0.00947f
C181 a_18_n7916# a_n33_n6777# 1.15e-19
C182 a_n76_5680# a_n76_6916# 0.00947f
C183 a_n76_n2972# a_18_n2972# 0.747f
C184 a_18_8152# w_n112_6816# 0.00199f
C185 a_n33_n1833# a_n33_n3069# 0.0665f
C186 a_n76_n9152# a_n33_n8013# 1.15e-19
C187 a_n33_n9249# a_n76_n7916# 1.15e-19
C188 w_n112_n5544# a_18_n4208# 0.00199f
C189 w_n112_n6780# a_n76_n7916# 0.00199f
C190 a_18_3208# a_n33_4347# 1.15e-19
C191 a_n33_8055# w_n112_6816# 4.13e-19
C192 w_n112_n5544# a_n76_n6680# 0.00199f
C193 a_n76_n9152# a_18_n9152# 0.747f
C194 a_n76_4444# w_n112_5580# 0.00199f
C195 a_n76_6916# w_n112_6816# 0.0182f
C196 a_18_1972# a_18_736# 0.00947f
C197 a_n33_639# a_n76_736# 0.0417f
C198 a_n76_n9152# w_n112_n10488# 0.00199f
C199 a_n33_n5541# a_n33_n6777# 0.0665f
C200 a_n33_n597# w_n112_n1836# 4.13e-19
C201 w_n112_4344# a_n33_3111# 4.13e-19
C202 a_18_n7916# w_n112_n9252# 0.00199f
C203 a_n33_n8013# a_n76_n7916# 0.0417f
C204 a_n76_n1736# w_n112_n600# 0.00199f
C205 a_n33_n597# w_n112_636# 4.13e-19
C206 a_18_n7916# a_18_n6680# 0.00947f
C207 a_n33_5583# a_n76_6916# 1.15e-19
C208 a_n76_n10388# w_n112_n9252# 0.00199f
C209 a_n76_n1736# a_n76_n2972# 0.00947f
C210 a_n33_n1833# a_18_n2972# 1.15e-19
C211 a_n33_4347# a_18_5680# 1.15e-19
C212 a_n76_5680# a_18_5680# 0.747f
C213 a_n33_n3069# a_n76_n4208# 1.15e-19
C214 a_n76_n2972# a_n33_n4305# 1.15e-19
C215 a_18_4444# w_n112_3108# 0.00199f
C216 a_18_n7916# a_n33_n9249# 1.15e-19
C217 w_n112_n6780# a_18_n7916# 0.00199f
C218 a_n76_n5444# a_n76_n6680# 0.00947f
C219 a_18_n5444# a_n33_n6777# 1.15e-19
C220 a_n33_n5541# a_18_n6680# 1.15e-19
C221 a_18_5680# w_n112_6816# 0.00199f
C222 a_n33_n9249# a_n76_n10388# 1.15e-19
C223 a_n76_n9152# a_n33_n10485# 1.15e-19
C224 a_n33_639# a_18_736# 0.0417f
C225 w_n112_n4308# a_n33_n3069# 4.13e-19
C226 a_n76_n500# w_n112_n1836# 0.00199f
C227 a_18_n1736# w_n112_n3072# 0.00199f
C228 a_18_9388# a_18_8152# 0.00947f
C229 w_n112_9288# a_n76_8152# 0.00199f
C230 a_n33_5583# a_18_5680# 0.0417f
C231 a_18_3208# w_n112_1872# 0.00199f
C232 a_18_n7916# a_n33_n8013# 0.0417f
C233 w_n112_n6780# a_n33_n5541# 4.13e-19
C234 a_n76_n500# w_n112_636# 0.00199f
C235 a_n33_n1833# a_n76_n1736# 0.0417f
C236 a_18_9388# a_n33_8055# 1.15e-19
C237 a_n33_n597# a_n76_n500# 0.0417f
C238 a_18_n7916# a_18_n9152# 0.00947f
C239 a_n76_9388# w_n112_9288# 0.0182f
C240 a_18_n5444# a_18_n6680# 0.00947f
C241 w_n112_3108# a_n33_4347# 4.13e-19
C242 a_n76_n10388# w_n112_n10488# 0.0182f
C243 w_n112_n4308# a_18_n2972# 0.00199f
C244 a_n76_4444# a_18_4444# 0.747f
C245 a_n76_736# a_18_736# 0.747f
C246 w_n112_n6780# a_18_n5444# 0.00199f
C247 a_18_n500# w_n112_n1836# 0.00199f
C248 a_n33_n3069# w_n112_n3072# 0.106f
C249 a_n33_8055# a_18_8152# 0.0417f
C250 a_n33_1875# w_n112_1872# 0.106f
C251 w_n112_n1836# a_n76_n2972# 0.00199f
C252 a_18_n500# w_n112_636# 0.00199f
C253 a_n33_n4305# a_n76_n4208# 0.0417f
C254 a_n33_n597# w_n112_n600# 0.106f
C255 w_n112_8052# a_n76_8152# 0.0182f
C256 a_n33_n597# a_18_n500# 0.0417f
C257 a_n33_8055# a_n76_6916# 1.15e-19
C258 w_n112_4344# a_18_4444# 0.0182f
C259 a_n76_3208# a_n33_4347# 1.15e-19
C260 a_n33_1875# w_n112_636# 4.13e-19
C261 a_n33_n6777# a_18_n6680# 0.0417f
C262 a_n33_n10485# a_n76_n10388# 0.0417f
C263 a_18_6916# w_n112_5580# 0.00199f
C264 a_n76_9388# w_n112_8052# 0.00199f
C265 w_n112_n5544# a_n76_n4208# 0.00199f
C266 w_n112_1872# a_n76_1972# 0.0182f
C267 w_n112_8052# a_18_6916# 0.00199f
C268 a_n76_4444# a_n76_5680# 0.00947f
C269 a_n76_4444# a_n33_4347# 0.0417f
C270 w_n112_n4308# a_n33_n4305# 0.106f
C271 a_n33_n5541# a_n33_n4305# 0.0665f
C272 a_18_n1736# a_n33_n3069# 1.15e-19
C273 a_n33_9291# w_n112_9288# 0.106f
C274 a_18_n2972# w_n112_n3072# 0.0182f
C275 a_n76_9388# a_n76_8152# 0.00947f
C276 w_n112_636# a_n76_1972# 0.00199f
C277 w_n112_n6780# a_n33_n6777# 0.106f
C278 a_n33_n1833# w_n112_n1836# 0.106f
C279 w_n112_n8016# a_n76_n6680# 0.00199f
C280 w_n112_n5544# a_n33_n5541# 0.106f
C281 a_18_4444# a_n33_3111# 1.15e-19
C282 w_n112_5580# a_n33_6819# 4.13e-19
C283 w_n112_8052# a_n33_6819# 4.13e-19
C284 a_n76_n500# w_n112_n600# 0.0182f
C285 a_n76_n500# a_18_n500# 0.747f
C286 a_n33_n597# a_n33_n1833# 0.0665f
C287 a_n76_n10388# a_18_n10388# 0.747f
C288 w_n112_4344# a_n76_5680# 0.00199f
C289 w_n112_4344# a_n33_4347# 0.106f
C290 a_n76_4444# a_n33_5583# 1.15e-19
C291 a_n33_n6777# a_n33_n8013# 0.0665f
C292 a_n76_n5444# a_n76_n4208# 0.00947f
C293 a_18_n5444# a_n33_n4305# 1.15e-19
C294 a_18_4444# w_n112_5580# 0.00199f
C295 a_n33_n9249# w_n112_n9252# 0.106f
C296 a_18_n1736# a_18_n2972# 0.00947f
C297 a_n76_8152# a_n33_6819# 1.15e-19
C298 w_n112_1872# a_18_1972# 0.0182f
C299 a_n76_n1736# w_n112_n3072# 0.00199f
C300 w_n112_n6780# a_18_n6680# 0.0182f
C301 a_n33_n4305# w_n112_n3072# 4.13e-19
C302 a_18_3208# a_n33_1875# 1.15e-19
C303 w_n112_n5544# a_18_n5444# 0.0182f
C304 a_n76_3208# w_n112_1872# 0.00199f
C305 w_n112_636# a_18_1972# 0.00199f
C306 a_n33_9291# w_n112_8052# 4.13e-19
C307 w_n112_n4308# a_n76_n5444# 0.00199f
C308 a_n33_n5541# a_n76_n5444# 0.0417f
C309 a_18_6916# a_n33_6819# 0.0417f
C310 a_18_n10388# VSUBS 0.426f
C311 a_n76_n10388# VSUBS 0.426f
C312 a_n33_n10485# VSUBS 0.192f
C313 a_18_n9152# VSUBS 0.415f
C314 a_n76_n9152# VSUBS 0.415f
C315 a_n33_n9249# VSUBS 0.156f
C316 a_18_n7916# VSUBS 0.415f
C317 a_n76_n7916# VSUBS 0.415f
C318 a_n33_n8013# VSUBS 0.156f
C319 a_18_n6680# VSUBS 0.415f
C320 a_n76_n6680# VSUBS 0.415f
C321 a_n33_n6777# VSUBS 0.156f
C322 a_18_n5444# VSUBS 0.415f
C323 a_n76_n5444# VSUBS 0.415f
C324 a_n33_n5541# VSUBS 0.156f
C325 a_18_n4208# VSUBS 0.415f
C326 a_n76_n4208# VSUBS 0.415f
C327 a_n33_n4305# VSUBS 0.156f
C328 a_18_n2972# VSUBS 0.415f
C329 a_n76_n2972# VSUBS 0.415f
C330 a_n33_n3069# VSUBS 0.156f
C331 a_18_n1736# VSUBS 0.415f
C332 a_n76_n1736# VSUBS 0.415f
C333 a_n33_n1833# VSUBS 0.156f
C334 a_18_n500# VSUBS 0.415f
C335 a_n76_n500# VSUBS 0.415f
C336 a_n33_n597# VSUBS 0.156f
C337 a_18_736# VSUBS 0.415f
C338 a_n76_736# VSUBS 0.415f
C339 a_n33_639# VSUBS 0.156f
C340 a_18_1972# VSUBS 0.415f
C341 a_n76_1972# VSUBS 0.415f
C342 a_n33_1875# VSUBS 0.156f
C343 a_18_3208# VSUBS 0.415f
C344 a_n76_3208# VSUBS 0.415f
C345 a_n33_3111# VSUBS 0.156f
C346 a_18_4444# VSUBS 0.415f
C347 a_n76_4444# VSUBS 0.415f
C348 a_n33_4347# VSUBS 0.156f
C349 a_18_5680# VSUBS 0.415f
C350 a_n76_5680# VSUBS 0.415f
C351 a_n33_5583# VSUBS 0.156f
C352 a_18_6916# VSUBS 0.415f
C353 a_n76_6916# VSUBS 0.415f
C354 a_n33_6819# VSUBS 0.156f
C355 a_18_8152# VSUBS 0.415f
C356 a_n76_8152# VSUBS 0.415f
C357 a_n33_8055# VSUBS 0.156f
C358 a_18_9388# VSUBS 0.426f
C359 a_n76_9388# VSUBS 0.426f
C360 a_n33_9291# VSUBS 0.192f
C361 w_n112_n10488# VSUBS 0.806f
C362 w_n112_n9252# VSUBS 0.806f
C363 w_n112_n8016# VSUBS 0.806f
C364 w_n112_n6780# VSUBS 0.806f
C365 w_n112_n5544# VSUBS 0.806f
C366 w_n112_n4308# VSUBS 0.806f
C367 w_n112_n3072# VSUBS 0.806f
C368 w_n112_n1836# VSUBS 0.806f
C369 w_n112_n600# VSUBS 0.806f
C370 w_n112_636# VSUBS 0.806f
C371 w_n112_1872# VSUBS 0.806f
C372 w_n112_3108# VSUBS 0.806f
C373 w_n112_4344# VSUBS 0.806f
C374 w_n112_5580# VSUBS 0.806f
C375 w_n112_6816# VSUBS 0.806f
C376 w_n112_8052# VSUBS 0.806f
C377 w_n112_9288# VSUBS 0.806f
.ends

.subckt sky130_fd_pr__pfet_01v8_F76D73 a_n1558_11242# a_n1558_n14714# a_n1500_n43239#
+ w_n1594_n3690# a_n1500_n11103# a_n1558_50794# a_1500_n23366# a_n1500_n50655# w_n1594_n56838#
+ w_n1594_n24702# a_1500_n30782# a_n1500_3729# a_n1558_n60446# w_n1594_12378# a_1500_n8534#
+ a_n1558_14950# a_1500_n19658# a_n1500_n14811# a_n1500_n46947# w_n1594_9906# w_n1594_n6162#
+ a_1500_22366# a_n1500_22269# a_n1558_53266# a_n1558_n56738# a_n1558_n24602# a_n1558_21130#
+ a_n1500_n53127# w_n1594_n13578# a_n1558_60682# a_1500_n33254# a_n1500_n60543# w_n1594_n20994#
+ a_1500_n40670# a_1500_18658# a_n1558_49558# a_n1558_17422# w_n1594_22266# a_n1500_n49419#
+ w_n1594_n9870# a_n1500_25977# a_n1558_56974# a_n1500_n56835# a_1500_n29546# a_n1558_n3590#
+ a_1500_n36962# a_n1500_9909# a_n1558_n13478# a_1500_32254# a_n1500_32157# a_n1558_n20894#
+ w_n1594_18558# w_n1594_n23466# a_1500_n43142# w_n1594_n30882# w_n1594_25974# a_n1500_n2451#
+ a_1500_28546# a_1500_n7298# a_n1500_28449# a_n1558_59446# a_n1558_27310# a_n1500_n13575#
+ a_n1500_n59307# w_n1594_32154# w_n1594_n19758# a_1500_35962# a_n1558_n6062# a_n1500_35865#
+ a_1500_n39434# a_n1500_n20991# a_1500_n46850# a_n1558_n23366# a_1500_42142# a_n1500_42045#
+ a_n1558_n30782# w_n1594_n33354# w_n1594_28446# a_1500_n53030# w_n1594_35862# w_n1594_n40770#
+ a_n1558_n9770# w_n1594_18# a_n1558_16186# a_n1500_21# a_n1558_n19658# a_n1500_n16047#
+ a_1500_38434# a_n1500_38337# a_n1500_n55599# a_n1500_n23463# w_n1594_n29646# a_1500_45850#
+ w_n1594_42042# a_n1500_45753# a_n1558_40906# a_1500_n49322# a_n1558_n33254# a_1500_52030#
+ a_n1500_n8631# a_n1558_n40670# a_n1558_19894# w_n1594_38334# w_n1594_n43242# a_n1500_n19755#
+ w_n1594_45750# a_n1558_26074# a_n1558_n29546# a_1500_48322# a_n1500_48225# a_1500_n38198#
+ a_n1558_33490# a_n1558_n36962# a_n1500_n33351# w_n1594_n39534# a_n1500_55641# a_1500_n59210#
+ w_n1594_n46950# a_n1558_n43142# a_n1558_29782# w_n1594_n53130# a_n1500_n29643# w_n1594_48222#
+ a_1500_37198# a_n1558_n39434# a_1500_58210# a_n1500_58113# a_n1500_12381# a_1500_n1118#
+ a_1500_n48086# a_n1558_n46850# w_n1594_n49422# a_n1500_n7395# a_n1558_n53030# w_n1594_37098#
+ a_n1558_39670# a_n1500_n39531# w_n1594_58110# a_1500_n4826# a_1500_47086# a_n1558_10006#
+ a_n1558_n49322# w_n1594_n2454# w_n1594_n38298# a_1500_2590# w_n1594_2490# w_n1594_n59310#
+ a_n1500_6201# a_n1500_18561# a_n1558_13714# a_n1558_2590# a_1500_n25838# a_n1558_n38198#
+ a_1500_5062# a_1500_118# a_n1558_n59210# w_n1594_n48186# w_n1594_n16050# a_1500_n32018#
+ a_n1500_2493# a_1500_24838# a_n1558_5062# a_n1500_n38295# w_n1594_n8634# a_1500_8770#
+ a_n1558_55738# a_n1558_23602# a_n1558_n2354# w_n1594_8670# a_1500_n35726# a_n1558_n48086#
+ a_1500_31018# w_n1594_n58074# w_n1594_24738# a_n1558_8770# a_n1500_n1215# a_n1558_12478#
+ a_n1500_n12339# a_n1500_n48183# a_1500_34726# a_n1500_34629# w_n1594_n25938# a_1500_n45614#
+ a_n1500_8673# w_n1594_n32118# a_n1500_n4923# w_n1594_34626# a_n1558_n8534# w_n1594_n7398#
+ a_n1558_22366# a_n1558_n25838# a_n1500_n22227# a_n1500_n58071# a_1500_44614# a_n1500_44517#
+ a_n1500_n61779# w_n1594_n35826# a_n1500_51933# a_1500_n55502# a_n1558_n32018# a_n1558_18658#
+ w_n1594_n42006# a_n1500_n18519# a_n1500_n25935# w_n1594_44514# w_n1594_51930# a_n1558_32254#
+ a_n1558_n35726# a_n1500_n32115# a_1500_54502# a_n1500_54405# a_1500_n44378# a_1500_n12242#
+ w_n1594_n45714# a_1500_n51794# a_n1500_n3687# a_n1558_28546# a_n1558_n7298# a_n1500_n28407#
+ a_n1558_35962# a_n1500_n35823# w_n1594_54402# a_1500_n15950# a_1500_43378# a_1500_11242#
+ a_n1500_11145# a_n1558_42142# a_n1558_n45614# a_1500_50794# a_n1500_n42003# a_n1500_50697#
+ a_1500_n54266# a_1500_n22130# a_n1500_n6159# w_n1594_n55602# a_1500_n61682# a_n1558_38434#
+ a_n1500_n24699# w_n1594_43278# w_n1594_11142# a_1500_14950# a_n1500_46989# a_n1558_45850#
+ a_n1500_14853# a_1500_n18422# a_n1500_n45711# w_n1594_50694# a_1500_n57974# a_n1500_n9867#
+ w_n1594_n1218# a_1500_53266# a_1500_1354# a_n1500_53169# a_1500_21130# a_n1500_21033#
+ a_n1558_n55502# a_n1558_52030# w_n1594_1254# w_n1594_n12342# w_n1594_n44478# a_1500_60682#
+ a_n1500_60585# w_n1594_14850# w_n1594_n51894# w_n1594_46986# a_1500_49558# a_1500_17422#
+ a_n1558_48322# a_n1500_17325# a_n1500_n34587# a_1500_56974# a_n1558_1354# w_n1594_53166#
+ w_n1594_21030# w_n1594_n4926# a_n1500_56877# a_n1500_24741# a_1500_n3590# a_1500_n28310#
+ w_n1594_60582# w_n1594_4962# a_n1558_n44378# a_n1558_n12242# a_n1558_n51794# w_n1594_17322#
+ w_n1594_n22230# w_n1594_n54366# w_n1594_49458# a_n1500_1257# w_n1594_n61782# w_n1594_56874#
+ a_n1558_37198# a_n1500_n37059# a_1500_59446# a_1500_27310# a_1500_7534# a_n1500_59349#
+ a_n1500_27213# a_1500_n6062# a_1500_n17186# a_n1558_58210# a_n1558_n15950# a_n1500_n44475#
+ a_n1558_n1118# w_n1594_7434# w_n1594_n18522# a_n1500_n51891# a_n1558_n54266# a_1500_n41906#
+ a_n1500_4965# a_n1558_n22130# a_n1558_n61682# w_n1594_59346# w_n1594_27210# a_n1558_7534#
+ a_1500_n9770# w_n1594_30918# a_n1558_n4826# a_1500_16186# a_n1500_16089# a_n1558_47086#
+ a_n1558_n18422# a_n1500_37101# a_n1558_n57974# a_1500_n27074# a_n1500_n54363# a_1500_40906#
+ w_n1594_n28410# a_n1500_40809# a_1500_n34490# a_n1500_7437# w_n1594_16086# a_1500_19894#
+ a_n1500_19797# w_n1594_40806# a_1500_26074# a_1500_6298# a_n1558_n28310# w_n1594_6198#
+ w_n1594_n17286# a_1500_33490# a_n1500_33393# w_n1594_19794# a_n1558_6298# a_1500_29782#
+ a_n1500_29685# a_n1558_24838# w_n1594_33390# a_n1558_n17186# a_n1558_118# a_n1558_31018#
+ w_n1594_n27174# a_n1500_43281# a_n1558_n41906# a_1500_n11006# w_n1594_29682# w_n1594_n34590#
+ a_1500_n50558# a_n1500_n17283# a_1500_39670# a_n1500_39573# a_n1558_34726# a_1500_n14714#
+ a_n1558_n27074# a_1500_10006# a_n1558_n34490# w_n1594_n37062# w_n1594_39570# a_1500_n60446#
+ a_n1500_n27171# a_1500_13714# a_n1500_13617# a_n1500_49461# a_n1558_44614# a_n1500_n30879#
+ a_1500_n56738# a_1500_n24602# w_n1594_n11106# w_n1594_n50658# w_n1594_13614# a_1500_55738#
+ a_1500_23602# a_1500_3826# a_n1500_23505# a_1500_n2354# a_1500_n13478# a_n1558_54502#
+ a_n1500_n40767# w_n1594_3726# w_n1594_n14814# a_n1500_30921# a_1500_n20894# a_n1558_n11006#
+ a_n1558_n50558# w_n1594_n60546# a_n1558_3826# w_n1594_55638# w_n1594_23502# VSUBS
+ a_1500_12478# a_n1558_43378#
X0 a_1500_53266# a_n1500_53169# a_n1558_53266# w_n1594_53166# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1 a_1500_n18422# a_n1500_n18519# a_n1558_n18422# w_n1594_n18522# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X2 a_1500_n45614# a_n1500_n45711# a_n1558_n45614# w_n1594_n45714# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X3 a_1500_n43142# a_n1500_n43239# a_n1558_n43142# w_n1594_n43242# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X4 a_1500_n22130# a_n1500_n22227# a_n1558_n22130# w_n1594_n22230# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X5 a_1500_n3590# a_n1500_n3687# a_n1558_n3590# w_n1594_n3690# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X6 a_1500_35962# a_n1500_35865# a_n1558_35962# w_n1594_35862# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X7 a_1500_33490# a_n1500_33393# a_n1558_33490# w_n1594_33390# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X8 a_1500_60682# a_n1500_60585# a_n1558_60682# w_n1594_60582# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X9 a_1500_12478# a_n1500_12381# a_n1558_12478# w_n1594_12378# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X10 a_1500_38434# a_n1500_38337# a_n1558_38434# w_n1594_38334# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X11 a_1500_6298# a_n1500_6201# a_n1558_6298# w_n1594_6198# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X12 a_1500_n55502# a_n1500_n55599# a_n1558_n55502# w_n1594_n55602# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X13 a_1500_n32018# a_n1500_n32115# a_n1558_n32018# w_n1594_n32118# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X14 a_1500_45850# a_n1500_45753# a_n1558_45850# w_n1594_45750# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X15 a_1500_24838# a_n1500_24741# a_n1558_24838# w_n1594_24738# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X16 a_1500_n38198# a_n1500_n38295# a_n1558_n38198# w_n1594_n38298# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X17 a_1500_22366# a_n1500_22269# a_n1558_22366# w_n1594_22266# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X18 a_1500_48322# a_n1500_48225# a_n1558_48322# w_n1594_48222# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X19 a_1500_n14714# a_n1500_n14811# a_n1558_n14714# w_n1594_n14814# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X20 a_1500_n41906# a_n1500_n42003# a_n1558_n41906# w_n1594_n42006# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X21 a_1500_n12242# a_n1500_n12339# a_n1558_n12242# w_n1594_n12342# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X22 a_1500_34726# a_n1500_34629# a_n1558_34726# w_n1594_34626# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X23 a_1500_32254# a_n1500_32157# a_n1558_32254# w_n1594_32154# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X24 a_1500_n48086# a_n1500_n48183# a_n1558_n48086# w_n1594_n48186# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X25 a_1500_58210# a_n1500_58113# a_n1558_58210# w_n1594_58110# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X26 a_1500_n24602# a_n1500_n24699# a_n1558_n24602# w_n1594_n24702# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X27 a_1500_14950# a_n1500_14853# a_n1558_14950# w_n1594_14850# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X28 a_1500_n8534# a_n1500_n8631# a_n1558_n8534# w_n1594_n8634# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X29 a_1500_n57974# a_n1500_n58071# a_n1558_n57974# w_n1594_n58074# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X30 a_1500_n6062# a_n1500_n6159# a_n1558_n6062# w_n1594_n6162# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X31 a_1500_n34490# a_n1500_n34587# a_n1558_n34490# w_n1594_n34590# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X32 a_1500_17422# a_n1500_17325# a_n1558_17422# w_n1594_17322# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X33 a_1500_44614# a_n1500_44517# a_n1558_44614# w_n1594_44514# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X34 a_1500_42142# a_n1500_42045# a_n1558_42142# w_n1594_42042# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X35 a_1500_8770# a_n1500_8673# a_n1558_8770# w_n1594_8670# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X36 a_1500_n11006# a_n1500_n11103# a_n1558_n11006# w_n1594_n11106# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X37 a_1500_n19658# a_n1500_n19755# a_n1558_n19658# w_n1594_n19758# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X38 a_1500_n46850# a_n1500_n46947# a_n1558_n46850# w_n1594_n46950# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X39 a_1500_n17186# a_n1500_n17283# a_n1558_n17186# w_n1594_n17286# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X40 a_1500_27310# a_n1500_27213# a_n1558_27310# w_n1594_27210# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X41 a_1500_n44378# a_n1500_n44475# a_n1558_n44378# w_n1594_n44478# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X42 a_1500_54502# a_n1500_54405# a_n1558_54502# w_n1594_54402# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X43 a_1500_52030# a_n1500_51933# a_n1558_52030# w_n1594_51930# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X44 a_1500_31018# a_n1500_30921# a_n1558_31018# w_n1594_30918# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X45 a_1500_n4826# a_n1500_n4923# a_n1558_n4826# w_n1594_n4926# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X46 a_1500_37198# a_n1500_37101# a_n1558_37198# w_n1594_37098# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X47 a_1500_n2354# a_n1500_n2451# a_n1558_n2354# w_n1594_n2454# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X48 a_1500_n51794# a_n1500_n51891# a_n1558_n51794# w_n1594_n51894# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X49 a_1500_n29546# a_n1500_n29643# a_n1558_n29546# w_n1594_n29646# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X50 a_1500_13714# a_n1500_13617# a_n1558_13714# w_n1594_13614# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X51 a_1500_n56738# a_n1500_n56835# a_n1558_n56738# w_n1594_n56838# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X52 a_1500_11242# a_n1500_11145# a_n1558_11242# w_n1594_11142# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X53 a_1500_40906# a_n1500_40809# a_n1558_40906# w_n1594_40806# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X54 a_1500_n27074# a_n1500_n27171# a_n1558_n27074# w_n1594_n27174# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X55 a_1500_n54266# a_n1500_n54363# a_n1558_n54266# w_n1594_n54366# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X56 a_1500_19894# a_n1500_19797# a_n1558_19894# w_n1594_19794# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X57 a_1500_2590# a_n1500_2493# a_n1558_2590# w_n1594_2490# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X58 a_1500_n59210# a_n1500_n59307# a_n1558_n59210# w_n1594_n59310# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X59 a_1500_7534# a_n1500_7437# a_n1558_7534# w_n1594_7434# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X60 a_1500_49558# a_n1500_49461# a_n1558_49558# w_n1594_49458# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X61 a_1500_n36962# a_n1500_n37059# a_n1558_n36962# w_n1594_n37062# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X62 a_1500_5062# a_n1500_4965# a_n1558_5062# w_n1594_4962# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X63 a_1500_47086# a_n1500_46989# a_n1558_47086# w_n1594_46986# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X64 a_1500_n15950# a_n1500_n16047# a_n1558_n15950# w_n1594_n16050# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X65 a_1500_n61682# a_n1500_n61779# a_n1558_n61682# w_n1594_n61782# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X66 a_1500_n13478# a_n1500_n13575# a_n1558_n13478# w_n1594_n13578# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X67 a_1500_23602# a_n1500_23505# a_n1558_23602# w_n1594_23502# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X68 a_1500_n40670# a_n1500_n40767# a_n1558_n40670# w_n1594_n40770# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X69 a_1500_n39434# a_n1500_n39531# a_n1558_n39434# w_n1594_n39534# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X70 a_1500_21130# a_n1500_21033# a_n1558_21130# w_n1594_21030# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X71 a_1500_29782# a_n1500_29685# a_n1558_29782# w_n1594_29682# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X72 a_1500_56974# a_n1500_56877# a_n1558_56974# w_n1594_56874# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X73 a_1500_59446# a_n1500_59349# a_n1558_59446# w_n1594_59346# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X74 a_1500_n20894# a_n1500_n20991# a_n1558_n20894# w_n1594_n20994# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X75 a_1500_n25838# a_n1500_n25935# a_n1558_n25838# w_n1594_n25938# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X76 a_1500_n23366# a_n1500_n23463# a_n1558_n23366# w_n1594_n23466# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X77 a_1500_n50558# a_n1500_n50655# a_n1558_n50558# w_n1594_n50658# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X78 a_1500_n49322# a_n1500_n49419# a_n1558_n49322# w_n1594_n49422# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X79 a_1500_n1118# a_n1500_n1215# a_n1558_n1118# w_n1594_n1218# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X80 a_1500_n9770# a_n1500_n9867# a_n1558_n9770# w_n1594_n9870# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X81 a_1500_n28310# a_n1500_n28407# a_n1558_n28310# w_n1594_n28410# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X82 a_1500_n7298# a_n1500_n7395# a_n1558_n7298# w_n1594_n7398# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X83 a_1500_10006# a_n1500_9909# a_n1558_10006# w_n1594_9906# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X84 a_1500_39670# a_n1500_39573# a_n1558_39670# w_n1594_39570# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X85 a_1500_18658# a_n1500_18561# a_n1558_18658# w_n1594_18558# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X86 a_1500_n53030# a_n1500_n53127# a_n1558_n53030# w_n1594_n53130# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X87 a_1500_3826# a_n1500_3729# a_n1558_3826# w_n1594_3726# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X88 a_1500_16186# a_n1500_16089# a_n1558_16186# w_n1594_16086# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X89 a_1500_1354# a_n1500_1257# a_n1558_1354# w_n1594_1254# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X90 a_1500_43378# a_n1500_43281# a_n1558_43378# w_n1594_43278# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X91 a_1500_n30782# a_n1500_n30879# a_n1558_n30782# w_n1594_n30882# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X92 a_1500_118# a_n1500_21# a_n1558_118# w_n1594_18# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X93 a_1500_n35726# a_n1500_n35823# a_n1558_n35726# w_n1594_n35826# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X94 a_1500_n33254# a_n1500_n33351# a_n1558_n33254# w_n1594_n33354# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X95 a_1500_n60446# a_n1500_n60543# a_n1558_n60446# w_n1594_n60546# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X96 a_1500_50794# a_n1500_50697# a_n1558_50794# w_n1594_50694# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X97 a_1500_28546# a_n1500_28449# a_n1558_28546# w_n1594_28446# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X98 a_1500_55738# a_n1500_55641# a_n1558_55738# w_n1594_55638# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X99 a_1500_26074# a_n1500_25977# a_n1558_26074# w_n1594_25974# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
C0 w_n1594_n22230# a_1500_n22130# 0.0187f
C1 a_n1500_44517# a_1500_44614# 0.217f
C2 a_n1500_n22227# a_1500_n22130# 0.217f
C3 w_n1594_2490# a_n1500_1257# 0.0172f
C4 a_n1500_n56835# a_n1500_n58071# 3.11f
C5 a_n1500_43281# w_n1594_43278# 1.65f
C6 a_1500_n36962# a_1500_n38198# 0.0105f
C7 a_n1500_n38295# a_n1558_n38198# 0.217f
C8 a_n1558_n41906# w_n1594_n43242# 0.0023f
C9 w_n1594_n54366# a_n1558_n53030# 0.0023f
C10 a_n1500_12381# w_n1594_12378# 1.65f
C11 w_n1594_39570# a_n1500_40809# 0.0172f
C12 a_n1500_38337# a_n1500_37101# 3.11f
C13 w_n1594_25974# a_n1500_24741# 0.0172f
C14 a_n1500_6201# w_n1594_6198# 1.65f
C15 a_n1500_n4923# a_1500_n4826# 0.217f
C16 a_n1500_n38295# w_n1594_n38298# 1.65f
C17 a_1500_55738# w_n1594_54402# 0.0023f
C18 a_n1500_54405# w_n1594_55638# 0.0172f
C19 a_n1500_n30879# a_n1500_n32115# 3.11f
C20 w_n1594_n61782# a_n1558_n60446# 0.0023f
C21 a_n1500_48225# a_n1558_48322# 0.217f
C22 w_n1594_n29646# a_n1558_n30782# 0.0023f
C23 a_n1558_n49322# w_n1594_n49422# 0.0187f
C24 w_n1594_n1218# a_n1558_n2354# 0.0023f
C25 a_n1500_55641# a_n1500_54405# 3.11f
C26 w_n1594_46986# a_1500_47086# 0.0187f
C27 w_n1594_22266# a_n1558_22366# 0.0187f
C28 w_n1594_n23466# a_n1558_n23366# 0.0187f
C29 a_n1558_32254# a_n1558_33490# 0.0105f
C30 a_n1500_n14811# w_n1594_n14814# 1.65f
C31 a_n1500_n11103# w_n1594_n11106# 1.65f
C32 a_n1558_n15950# w_n1594_n17286# 0.0023f
C33 a_1500_n53030# a_1500_n54266# 0.0105f
C34 a_n1500_n54363# a_n1558_n54266# 0.217f
C35 a_1500_n14714# a_1500_n15950# 0.0105f
C36 a_n1500_n16047# a_n1558_n15950# 0.217f
C37 a_n1558_n24602# a_n1558_n25838# 0.0105f
C38 a_n1500_30921# w_n1594_30918# 1.65f
C39 a_n1500_60585# a_1500_60682# 0.217f
C40 a_1500_5062# w_n1594_3726# 0.0023f
C41 a_n1558_3826# w_n1594_2490# 0.0023f
C42 a_n1558_42142# a_n1558_40906# 0.0105f
C43 w_n1594_35862# a_n1558_34726# 0.0023f
C44 w_n1594_34626# a_n1558_35962# 0.0023f
C45 w_n1594_51930# a_n1558_50794# 0.0023f
C46 a_n1558_n7298# a_n1558_n8534# 0.0105f
C47 a_1500_n39434# w_n1594_n40770# 0.0023f
C48 w_n1594_28446# a_n1500_28449# 1.65f
C49 a_1500_n13478# w_n1594_n13578# 0.0187f
C50 w_n1594_24738# a_n1500_24741# 1.65f
C51 a_n1500_4965# a_n1500_3729# 3.11f
C52 a_n1500_27213# a_n1558_27310# 0.217f
C53 a_1500_28546# a_1500_27310# 0.0105f
C54 a_n1558_42142# w_n1594_40806# 0.0023f
C55 a_n1500_19797# a_n1558_19894# 0.217f
C56 a_1500_21130# a_1500_19894# 0.0105f
C57 a_n1558_n18422# w_n1594_n18522# 0.0187f
C58 a_n1558_n35726# w_n1594_n35826# 0.0187f
C59 w_n1594_9906# a_n1558_11242# 0.0023f
C60 w_n1594_n27174# a_n1500_n28407# 0.0172f
C61 w_n1594_n59310# a_1500_n57974# 0.0023f
C62 w_n1594_25974# a_n1500_27213# 0.0172f
C63 w_n1594_n7398# a_1500_n7298# 0.0187f
C64 a_n1500_n48183# a_n1500_n49419# 3.11f
C65 a_n1500_n9867# a_n1500_n11103# 3.11f
C66 w_n1594_18558# a_n1500_18561# 1.65f
C67 a_n1500_n16047# w_n1594_n16050# 1.65f
C68 a_n1500_44517# w_n1594_45750# 0.0172f
C69 w_n1594_27210# a_1500_26074# 0.0023f
C70 a_1500_48322# a_1500_47086# 0.0105f
C71 a_1500_n46850# w_n1594_n46950# 0.0187f
C72 a_n1500_46989# a_n1558_47086# 0.217f
C73 a_1500_n44378# w_n1594_n45714# 0.0023f
C74 w_n1594_29682# a_n1500_28449# 0.0172f
C75 w_n1594_42042# a_1500_42142# 0.0187f
C76 w_n1594_n56838# a_1500_n55502# 0.0023f
C77 a_n1558_7534# w_n1594_8670# 0.0023f
C78 a_1500_n59210# a_1500_n60446# 0.0105f
C79 a_n1558_60682# w_n1594_59346# 0.0023f
C80 w_n1594_18# a_n1558_118# 0.0187f
C81 a_n1500_n60543# a_n1558_n60446# 0.217f
C82 a_1500_n1118# a_1500_n2354# 0.0105f
C83 w_n1594_23502# a_n1558_23602# 0.0187f
C84 a_n1500_n2451# a_n1558_n2354# 0.217f
C85 a_n1558_n20894# w_n1594_n20994# 0.0187f
C86 a_n1558_11242# a_n1558_10006# 0.0105f
C87 w_n1594_38334# a_1500_37198# 0.0023f
C88 a_n1558_10006# w_n1594_11142# 0.0023f
C89 a_n1500_n28407# a_1500_n28310# 0.217f
C90 a_n1500_n9867# w_n1594_n9870# 1.65f
C91 a_n1500_n44475# a_n1558_n44378# 0.217f
C92 a_1500_n51794# w_n1594_n51894# 0.0187f
C93 a_1500_n43142# a_1500_n44378# 0.0105f
C94 w_n1594_n30882# a_n1558_n29546# 0.0023f
C95 a_n1558_34726# w_n1594_33390# 0.0023f
C96 w_n1594_n33354# a_1500_n32018# 0.0023f
C97 a_n1558_6298# w_n1594_7434# 0.0023f
C98 w_n1594_19794# a_n1500_21033# 0.0172f
C99 a_n1558_48322# a_n1558_47086# 0.0105f
C100 a_1500_n33254# w_n1594_n33354# 0.0187f
C101 w_n1594_21030# a_1500_22366# 0.0023f
C102 w_n1594_n25938# a_n1500_n27171# 0.0172f
C103 w_n1594_2490# a_1500_1354# 0.0023f
C104 a_n1558_n56738# a_n1558_n57974# 0.0105f
C105 w_n1594_n22230# a_n1558_n23366# 0.0023f
C106 a_n1500_25977# a_n1500_24741# 3.11f
C107 a_1500_43378# w_n1594_43278# 0.0187f
C108 a_n1500_n38295# a_n1500_n39531# 3.11f
C109 a_n1500_n43239# w_n1594_n43242# 1.65f
C110 w_n1594_50694# a_n1500_51933# 0.0172f
C111 w_n1594_n54366# a_n1500_n54363# 1.65f
C112 a_n1558_38434# a_n1558_37198# 0.0105f
C113 a_1500_12478# w_n1594_12378# 0.0187f
C114 a_1500_6298# w_n1594_6198# 0.0187f
C115 a_1500_n38198# w_n1594_n38298# 0.0187f
C116 a_1500_54502# w_n1594_55638# 0.0023f
C117 a_n1558_54502# w_n1594_54402# 0.0187f
C118 a_n1500_7437# a_1500_7534# 0.217f
C119 w_n1594_14850# a_n1558_13714# 0.0023f
C120 a_n1558_58210# w_n1594_56874# 0.0023f
C121 a_n1500_58113# a_n1500_59349# 3.11f
C122 a_n1558_n30782# a_n1558_n32018# 0.0105f
C123 w_n1594_n61782# a_n1500_n61779# 1.65f
C124 a_n1500_24741# a_n1558_24838# 0.217f
C125 w_n1594_n28410# a_n1500_n27171# 0.0172f
C126 a_n1558_53266# w_n1594_54402# 0.0023f
C127 a_n1500_n50655# w_n1594_n49422# 0.0172f
C128 a_n1558_55738# a_n1558_54502# 0.0105f
C129 w_n1594_46986# a_n1558_45850# 0.0023f
C130 w_n1594_22266# a_n1500_21033# 0.0172f
C131 w_n1594_n23466# a_n1500_n24699# 0.0172f
C132 a_1500_n14714# w_n1594_n14814# 0.0187f
C133 a_1500_n11006# w_n1594_n11106# 0.0187f
C134 a_n1500_n17283# w_n1594_n17286# 1.65f
C135 a_n1500_n54363# a_n1500_n55599# 3.11f
C136 w_n1594_n3690# a_n1558_n2354# 0.0023f
C137 a_n1500_n16047# a_n1500_n17283# 3.11f
C138 a_1500_n24602# a_1500_n25838# 0.0105f
C139 a_n1500_n25935# a_n1558_n25838# 0.217f
C140 a_1500_31018# w_n1594_30918# 0.0187f
C141 a_n1500_40809# a_n1558_40906# 0.217f
C142 a_n1558_3826# w_n1594_3726# 0.0187f
C143 a_n1500_2493# w_n1594_2490# 1.65f
C144 a_1500_58210# w_n1594_59346# 0.0023f
C145 w_n1594_34626# a_n1500_34629# 1.65f
C146 a_n1500_34629# a_1500_34726# 0.217f
C147 a_n1500_n1215# w_n1594_n2454# 0.0172f
C148 a_1500_n7298# a_1500_n8534# 0.0105f
C149 w_n1594_28446# a_1500_28546# 0.0187f
C150 a_n1558_n40670# w_n1594_n40770# 0.0187f
C151 a_n1500_n8631# a_n1558_n8534# 0.217f
C152 a_n1558_n14714# w_n1594_n13578# 0.0023f
C153 a_n1558_5062# a_n1558_3826# 0.0105f
C154 a_n1500_27213# a_n1500_25977# 3.11f
C155 a_n1500_40809# w_n1594_40806# 1.65f
C156 a_n1500_19797# a_n1500_18561# 3.11f
C157 a_n1500_n19755# w_n1594_n18522# 0.0172f
C158 a_n1500_n37059# w_n1594_n35826# 0.0172f
C159 a_n1558_33490# w_n1594_32154# 0.0023f
C160 w_n1594_9906# a_n1500_9909# 1.65f
C161 w_n1594_n59310# a_n1558_n59210# 0.0187f
C162 w_n1594_n20994# a_1500_n20894# 0.0187f
C163 w_n1594_n27174# a_1500_n28310# 0.0023f
C164 w_n1594_25974# a_1500_27310# 0.0023f
C165 w_n1594_n7398# a_n1558_n8534# 0.0023f
C166 w_n1594_18558# a_1500_18658# 0.0187f
C167 a_n1558_n48086# a_n1558_n49322# 0.0105f
C168 a_1500_n15950# w_n1594_n16050# 0.0187f
C169 a_n1558_n9770# a_n1558_n11006# 0.0105f
C170 a_1500_44614# w_n1594_45750# 0.0023f
C171 a_n1500_46989# a_n1500_45753# 3.11f
C172 a_n1558_n48086# w_n1594_n46950# 0.0023f
C173 a_n1500_40809# a_1500_40906# 0.217f
C174 a_n1500_n35823# a_1500_n35726# 0.217f
C175 w_n1594_29682# a_1500_28546# 0.0023f
C176 w_n1594_n56838# a_n1558_n56738# 0.0187f
C177 w_n1594_42042# a_n1558_40906# 0.0023f
C178 a_n1500_n60543# a_n1500_n61779# 3.11f
C179 a_n1500_n2451# a_n1500_n3687# 3.11f
C180 w_n1594_23502# a_n1500_22269# 0.0172f
C181 a_1500_11242# a_1500_10006# 0.0105f
C182 w_n1594_n9870# a_n1500_n8631# 0.0172f
C183 a_n1500_9909# a_n1558_10006# 0.217f
C184 a_n1500_50697# a_1500_50794# 0.217f
C185 a_n1558_n11006# w_n1594_n12342# 0.0023f
C186 a_1500_n9770# w_n1594_n9870# 0.0187f
C187 w_n1594_n30882# a_n1500_n30879# 1.65f
C188 a_n1558_n53030# w_n1594_n51894# 0.0023f
C189 a_n1500_n49419# w_n1594_n50658# 0.0172f
C190 a_n1500_33393# w_n1594_33390# 1.65f
C191 a_n1500_n20991# a_n1500_n22227# 3.11f
C192 a_n1500_n20991# w_n1594_n22230# 0.0172f
C193 w_n1594_19794# a_1500_21130# 0.0023f
C194 a_n1558_n34490# w_n1594_n33354# 0.0023f
C195 w_n1594_42042# a_1500_40906# 0.0023f
C196 a_n1500_n51891# a_1500_n51794# 0.217f
C197 w_n1594_n56838# a_1500_n56738# 0.0187f
C198 a_n1500_n13575# a_1500_n13478# 0.217f
C199 w_n1594_21030# a_n1558_21130# 0.0187f
C200 w_n1594_n25938# a_1500_n27074# 0.0023f
C201 w_n1594_n24702# a_n1558_n23366# 0.0023f
C202 a_1500_n45614# w_n1594_n44478# 0.0023f
C203 a_n1558_42142# w_n1594_43278# 0.0023f
C204 a_1500_n43142# w_n1594_n43242# 0.0187f
C205 a_n1558_n38198# a_n1558_n39434# 0.0105f
C206 a_1500_38434# a_1500_37198# 0.0105f
C207 w_n1594_n54366# a_1500_n54266# 0.0187f
C208 a_n1558_13714# w_n1594_13614# 0.0187f
C209 w_n1594_50694# a_1500_52030# 0.0023f
C210 a_n1500_37101# a_n1558_37198# 0.217f
C211 a_n1558_11242# w_n1594_12378# 0.0023f
C212 a_n1558_5062# w_n1594_6198# 0.0023f
C213 a_n1500_39573# a_1500_39670# 0.217f
C214 a_n1558_n39434# w_n1594_n38298# 0.0023f
C215 a_n1500_n35823# w_n1594_n37062# 0.0172f
C216 a_n1500_29685# a_1500_29782# 0.217f
C217 a_1500_n30782# a_1500_n32018# 0.0105f
C218 w_n1594_n61782# a_1500_n61682# 0.0187f
C219 a_n1500_22269# a_1500_22366# 0.217f
C220 a_n1500_n32115# a_n1558_n32018# 0.217f
C221 a_n1500_24741# a_n1500_23505# 3.11f
C222 w_n1594_n28410# a_1500_n27074# 0.0023f
C223 a_n1500_n44475# a_n1500_n45711# 3.11f
C224 a_1500_n50558# w_n1594_n49422# 0.0023f
C225 a_1500_59446# w_n1594_59346# 0.0187f
C226 a_n1558_n46850# w_n1594_n48186# 0.0023f
C227 a_1500_55738# a_1500_54502# 0.0105f
C228 a_n1500_54405# a_n1558_54502# 0.217f
C229 w_n1594_22266# a_1500_21130# 0.0023f
C230 w_n1594_n1218# a_n1500_21# 0.0172f
C231 w_n1594_n23466# a_1500_n24602# 0.0023f
C232 a_1500_60682# w_n1594_60582# 0.0187f
C233 a_n1500_n58071# a_1500_n57974# 0.217f
C234 a_n1558_n15950# w_n1594_n14814# 0.0023f
C235 w_n1594_1254# a_n1500_1257# 1.65f
C236 a_n1558_n12242# w_n1594_n11106# 0.0023f
C237 a_1500_n17186# w_n1594_n17286# 0.0187f
C238 a_n1558_n54266# a_n1558_n55502# 0.0105f
C239 w_n1594_n3690# a_n1500_n3687# 1.65f
C240 a_n1558_n15950# a_n1558_n17186# 0.0105f
C241 w_n1594_14850# a_n1558_16186# 0.0023f
C242 a_n1500_n25935# a_n1500_n27171# 3.11f
C243 a_n1558_29782# w_n1594_30918# 0.0023f
C244 a_n1500_2493# w_n1594_3726# 0.0172f
C245 a_n1500_53169# a_n1558_53266# 0.217f
C246 a_n1558_n51794# w_n1594_n53130# 0.0023f
C247 a_n1500_56877# w_n1594_58110# 0.0172f
C248 a_n1500_n42003# a_1500_n41906# 0.217f
C249 w_n1594_34626# a_1500_34726# 0.0187f
C250 a_1500_n1118# w_n1594_n2454# 0.0023f
C251 a_n1500_n42003# w_n1594_n40770# 0.0172f
C252 w_n1594_28446# a_n1558_27310# 0.0023f
C253 a_n1500_n18519# w_n1594_n19758# 0.0172f
C254 a_1500_5062# a_1500_3826# 0.0105f
C255 a_n1500_3729# a_n1558_3826# 0.217f
C256 a_n1558_27310# a_n1558_26074# 0.0105f
C257 a_1500_n36962# w_n1594_n35826# 0.0023f
C258 a_n1558_19894# a_n1558_18658# 0.0105f
C259 a_1500_n19658# w_n1594_n18522# 0.0023f
C260 a_n1558_n33254# w_n1594_n34590# 0.0023f
C261 w_n1594_9906# a_1500_10006# 0.0187f
C262 w_n1594_n59310# a_n1500_n60543# 0.0172f
C263 w_n1594_25974# a_n1558_26074# 0.0187f
C264 w_n1594_17322# a_n1500_18561# 0.0172f
C265 w_n1594_18558# a_n1558_17422# 0.0023f
C266 a_n1500_n49419# a_n1558_n49322# 0.217f
C267 a_1500_n48086# a_1500_n49322# 0.0105f
C268 a_1500_n9770# a_1500_n11006# 0.0105f
C269 a_n1500_n11103# a_n1558_n11006# 0.217f
C270 a_n1558_n17186# w_n1594_n16050# 0.0023f
C271 a_n1558_47086# a_n1558_45850# 0.0105f
C272 w_n1594_44514# a_n1500_45753# 0.0172f
C273 a_n1500_58113# a_n1558_58210# 0.217f
C274 a_1500_59446# a_1500_58210# 0.0105f
C275 a_n1558_n60446# a_n1558_n61682# 0.0105f
C276 w_n1594_25974# a_1500_24838# 0.0023f
C277 w_n1594_23502# a_1500_22366# 0.0023f
C278 a_n1558_n2354# a_n1558_n3590# 0.0105f
C279 a_n1500_6201# w_n1594_4962# 0.0172f
C280 a_n1558_n38198# w_n1594_n39534# 0.0023f
C281 a_n1500_1257# a_n1558_1354# 0.217f
C282 a_1500_2590# a_1500_1354# 0.0105f
C283 a_n1500_n19755# a_1500_n19658# 0.217f
C284 w_n1594_n9870# a_1500_n8534# 0.0023f
C285 a_n1500_9909# a_n1500_8673# 3.11f
C286 a_n1500_32157# a_n1558_32254# 0.217f
C287 a_1500_33490# a_1500_32254# 0.0105f
C288 w_n1594_48222# a_n1500_49461# 0.0172f
C289 a_n1558_n11006# w_n1594_n9870# 0.0023f
C290 a_n1500_n12339# w_n1594_n12342# 1.65f
C291 w_n1594_n30882# a_1500_n30782# 0.0187f
C292 a_1500_n49322# w_n1594_n50658# 0.0023f
C293 a_n1558_n20894# a_n1558_n22130# 0.0105f
C294 w_n1594_19794# a_n1558_19894# 0.0187f
C295 a_n1500_16089# a_1500_16186# 0.217f
C296 w_n1594_39570# a_n1500_39573# 1.65f
C297 w_n1594_37098# a_n1500_38337# 0.0172f
C298 a_n1500_54405# w_n1594_53166# 0.0172f
C299 w_n1594_n56838# a_n1558_n57974# 0.0023f
C300 w_n1594_24738# a_n1558_26074# 0.0023f
C301 w_n1594_18# a_n1558_n1118# 0.0023f
C302 w_n1594_21030# a_n1500_19797# 0.0172f
C303 w_n1594_n6162# a_n1558_n4826# 0.0023f
C304 a_n1500_43281# a_1500_43378# 0.217f
C305 w_n1594_n24702# a_n1500_n24699# 1.65f
C306 a_n1500_53169# w_n1594_53166# 1.65f
C307 a_n1500_n23463# a_1500_n23366# 0.217f
C308 a_n1558_118# a_n1558_n1118# 0.0105f
C309 a_1500_n38198# a_1500_n39434# 0.0105f
C310 a_n1558_n44378# w_n1594_n43242# 0.0023f
C311 a_n1500_n39531# a_n1558_n39434# 0.217f
C312 w_n1594_49458# a_n1558_50794# 0.0023f
C313 a_n1500_n40767# w_n1594_n42006# 0.0172f
C314 a_n1500_37101# a_n1500_35865# 3.11f
C315 w_n1594_50694# a_n1558_50794# 0.0187f
C316 a_n1500_12381# w_n1594_13614# 0.0172f
C317 a_n1500_n6159# a_1500_n6062# 0.217f
C318 w_n1594_n54366# a_n1558_n55502# 0.0023f
C319 w_n1594_24738# a_1500_24838# 0.0187f
C320 a_n1500_2493# a_1500_2590# 0.217f
C321 a_1500_n35726# w_n1594_n37062# 0.0023f
C322 a_n1500_n7395# w_n1594_n8634# 0.0172f
C323 a_n1500_n32115# a_n1500_n33351# 3.11f
C324 w_n1594_n60546# a_n1500_n59307# 0.0172f
C325 w_n1594_n28410# a_n1558_n28310# 0.0187f
C326 a_n1500_n48183# w_n1594_n48186# 1.65f
C327 w_n1594_n58074# a_n1500_n56835# 0.0172f
C328 w_n1594_n4926# a_n1500_n3687# 0.0172f
C329 w_n1594_1254# a_1500_1354# 0.0187f
C330 a_1500_n54266# a_1500_n55502# 0.0105f
C331 a_n1500_n55599# a_n1558_n55502# 0.217f
C332 a_n1558_n18422# w_n1594_n17286# 0.0023f
C333 a_1500_n15950# a_1500_n17186# 0.0105f
C334 a_n1500_12381# a_1500_12478# 0.217f
C335 w_n1594_n3690# a_1500_n3590# 0.0187f
C336 a_n1500_n17283# a_n1558_n17186# 0.217f
C337 w_n1594_14850# a_n1500_14853# 1.65f
C338 a_n1558_n25838# a_n1558_n27074# 0.0105f
C339 a_n1500_53169# a_n1500_51933# 3.11f
C340 a_1500_56974# w_n1594_58110# 0.0023f
C341 a_n1500_n53127# w_n1594_n53130# 1.65f
C342 w_n1594_34626# a_n1558_33490# 0.0023f
C343 w_n1594_16086# a_n1500_17325# 0.0172f
C344 a_n1558_n2354# w_n1594_n2454# 0.0187f
C345 a_1500_n41906# w_n1594_n40770# 0.0023f
C346 w_n1594_n34590# a_n1500_n33351# 0.0172f
C347 a_1500_n18422# w_n1594_n19758# 0.0023f
C348 a_n1500_3729# a_n1500_2493# 3.11f
C349 a_n1500_25977# a_n1558_26074# 0.217f
C350 a_1500_27310# a_1500_26074# 0.0105f
C351 a_1500_19894# a_1500_18658# 0.0105f
C352 a_n1500_18561# a_n1558_18658# 0.217f
C353 a_n1500_n34587# w_n1594_n34590# 1.65f
C354 w_n1594_n1218# a_n1558_118# 0.0023f
C355 w_n1594_n59310# a_1500_n60446# 0.0023f
C356 w_n1594_9906# a_n1558_8770# 0.0023f
C357 a_n1500_n49419# a_n1500_n50655# 3.11f
C358 w_n1594_17322# a_1500_18658# 0.0023f
C359 a_n1500_n11103# a_n1500_n12339# 3.11f
C360 a_1500_47086# a_1500_45850# 0.0105f
C361 a_n1500_45753# a_n1558_45850# 0.217f
C362 a_n1558_26074# a_n1558_24838# 0.0105f
C363 a_n1558_n45614# w_n1594_n45714# 0.0187f
C364 a_n1500_n45711# w_n1594_n46950# 0.0172f
C365 w_n1594_44514# a_1500_45850# 0.0023f
C366 a_n1558_n43142# w_n1594_n44478# 0.0023f
C367 a_1500_n60446# a_1500_n61682# 0.0105f
C368 w_n1594_n55602# a_n1558_n54266# 0.0023f
C369 a_n1500_n61779# a_n1558_n61682# 0.217f
C370 a_1500_n2354# a_1500_n3590# 0.0105f
C371 a_n1500_2493# w_n1594_1254# 0.0172f
C372 a_n1500_n3687# a_n1558_n3590# 0.217f
C373 a_n1500_56877# w_n1594_56874# 1.65f
C374 a_n1500_n39531# w_n1594_n39534# 1.65f
C375 a_1500_6298# w_n1594_4962# 0.0023f
C376 a_n1500_1257# a_n1500_21# 3.11f
C377 a_n1558_10006# a_n1558_8770# 0.0105f
C378 a_n1500_32157# a_n1500_30921# 3.11f
C379 a_n1500_n29643# a_1500_n29546# 0.217f
C380 w_n1594_48222# a_1500_49558# 0.0023f
C381 a_n1500_59349# a_n1558_59446# 0.217f
C382 a_1500_n12242# w_n1594_n12342# 0.0187f
C383 w_n1594_n30882# a_n1558_n32018# 0.0023f
C384 w_n1594_n29646# a_n1500_n28407# 0.0172f
C385 a_n1558_n50558# w_n1594_n50658# 0.0187f
C386 a_n1500_56877# a_1500_56974# 0.217f
C387 w_n1594_19794# a_n1500_18561# 0.0172f
C388 a_1500_54502# w_n1594_53166# 0.0023f
C389 w_n1594_37098# a_1500_38434# 0.0023f
C390 w_n1594_21030# a_1500_19894# 0.0023f
C391 w_n1594_n24702# a_1500_n24602# 0.0187f
C392 w_n1594_n6162# a_n1500_n6159# 1.65f
C393 a_n1500_32157# w_n1594_32154# 1.65f
C394 a_1500_53266# w_n1594_53166# 0.0187f
C395 a_1500_118# a_1500_n1118# 0.0105f
C396 a_n1500_n39531# a_n1500_n40767# 3.11f
C397 w_n1594_35862# a_n1500_37101# 0.0172f
C398 a_1500_n40670# w_n1594_n42006# 0.0023f
C399 a_n1558_37198# a_n1558_35962# 0.0105f
C400 w_n1594_49458# a_n1500_49461# 1.65f
C401 w_n1594_50694# a_n1500_49461# 0.0172f
C402 a_1500_12478# w_n1594_13614# 0.0023f
C403 w_n1594_51930# a_n1500_53169# 0.0172f
C404 w_n1594_24738# a_n1558_23602# 0.0023f
C405 a_n1500_6201# a_1500_6298# 0.217f
C406 a_n1558_n36962# w_n1594_n37062# 0.0187f
C407 a_1500_n7298# w_n1594_n8634# 0.0023f
C408 w_n1594_n60546# a_1500_n59210# 0.0023f
C409 w_n1594_n28410# a_n1500_n29643# 0.0172f
C410 a_n1500_n46947# a_1500_n46850# 0.217f
C411 a_n1558_n9770# w_n1594_n8634# 0.0023f
C412 a_1500_n33254# a_n1500_n33351# 0.217f
C413 w_n1594_27210# a_n1558_28546# 0.0023f
C414 a_1500_n48086# w_n1594_n48186# 0.0187f
C415 a_1500_33490# w_n1594_33390# 0.0187f
C416 a_n1558_n33254# a_n1558_n34490# 0.0105f
C417 a_n1500_9909# w_n1594_8670# 0.0172f
C418 w_n1594_n4926# a_1500_n3590# 0.0023f
C419 a_n1500_n55599# a_n1500_n56835# 3.11f
C420 w_n1594_13614# a_n1500_14853# 0.0172f
C421 a_n1500_n17283# a_n1500_n18519# 3.11f
C422 a_n1500_39573# w_n1594_40806# 0.0172f
C423 w_n1594_n3690# a_n1558_n4826# 0.0023f
C424 w_n1594_38334# a_n1558_39670# 0.0023f
C425 a_n1500_12381# w_n1594_11142# 0.0172f
C426 w_n1594_14850# a_1500_14950# 0.0187f
C427 a_n1500_n27171# a_n1558_n27074# 0.217f
C428 a_1500_n25838# a_1500_n27074# 0.0105f
C429 a_n1558_53266# a_n1558_52030# 0.0105f
C430 w_n1594_n32118# a_n1558_n30782# 0.0023f
C431 a_1500_n53030# w_n1594_n53130# 0.0187f
C432 w_n1594_16086# a_1500_17422# 0.0023f
C433 a_n1500_n3687# w_n1594_n2454# 0.0172f
C434 w_n1594_n20994# a_n1500_n22227# 0.0172f
C435 a_n1558_n19658# w_n1594_n19758# 0.0187f
C436 a_n1500_8673# w_n1594_7434# 0.0172f
C437 w_n1594_48222# a_n1500_46989# 0.0172f
C438 a_n1558_3826# a_n1558_2590# 0.0105f
C439 a_n1500_18561# a_n1500_17325# 3.11f
C440 a_1500_n34490# w_n1594_n34590# 0.0187f
C441 w_n1594_n58074# a_n1500_n58071# 1.65f
C442 a_n1558_n49322# a_n1558_n50558# 0.0105f
C443 w_n1594_17322# a_n1558_17422# 0.0187f
C444 a_n1558_n11006# a_n1558_n12242# 0.0105f
C445 a_1500_26074# a_1500_24838# 0.0105f
C446 a_n1500_45753# a_n1500_44517# 3.11f
C447 a_1500_13714# a_n1500_13617# 0.217f
C448 a_n1500_n46947# w_n1594_n45714# 0.0172f
C449 w_n1594_44514# a_n1558_44614# 0.0187f
C450 a_n1500_n37059# a_1500_n36962# 0.217f
C451 a_n1500_n44475# w_n1594_n44478# 1.65f
C452 w_n1594_n55602# a_n1500_n55599# 1.65f
C453 a_n1500_n3687# a_n1500_n4923# 3.11f
C454 a_n1558_5062# w_n1594_4962# 0.0187f
C455 a_1500_n39434# w_n1594_n39534# 0.0187f
C456 a_n1558_56974# w_n1594_55638# 0.0023f
C457 a_1500_56974# w_n1594_56874# 0.0187f
C458 a_1500_10006# a_1500_8770# 0.0105f
C459 a_n1558_32254# a_n1558_31018# 0.0105f
C460 a_n1500_8673# a_n1558_8770# 0.217f
C461 a_n1558_24838# a_n1558_23602# 0.0105f
C462 w_n1594_48222# a_n1558_48322# 0.0187f
C463 a_n1500_49461# a_1500_49558# 0.217f
C464 a_n1558_n13478# w_n1594_n12342# 0.0023f
C465 a_n1558_n44378# a_n1558_n45614# 0.0105f
C466 a_n1500_n51891# w_n1594_n50658# 0.0172f
C467 a_n1500_58113# w_n1594_58110# 1.65f
C468 w_n1594_n29646# a_1500_n28310# 0.0023f
C469 w_n1594_19794# a_1500_18658# 0.0023f
C470 a_n1500_59349# w_n1594_59346# 1.65f
C471 w_n1594_37098# a_n1558_37198# 0.0187f
C472 a_n1500_n53127# a_1500_n53030# 0.217f
C473 a_n1500_n14811# a_1500_n14714# 0.217f
C474 a_1500_32254# w_n1594_32154# 0.0187f
C475 w_n1594_n6162# a_1500_n6062# 0.0187f
C476 w_n1594_18# a_n1500_1257# 0.0172f
C477 w_n1594_n24702# a_n1558_n25838# 0.0023f
C478 a_n1558_52030# w_n1594_53166# 0.0023f
C479 w_n1594_35862# a_1500_37198# 0.0023f
C480 a_n1558_n39434# a_n1558_n40670# 0.0105f
C481 a_n1558_n41906# w_n1594_n42006# 0.0187f
C482 a_1500_37198# a_1500_35962# 0.0105f
C483 a_n1500_35865# a_n1558_35962# 0.217f
C484 w_n1594_49458# a_1500_49558# 0.0187f
C485 w_n1594_50694# a_1500_49558# 0.0023f
C486 w_n1594_51930# a_1500_53266# 0.0023f
C487 a_n1500_n12339# w_n1594_n13578# 0.0172f
C488 a_n1500_n38295# w_n1594_n37062# 0.0172f
C489 a_n1500_28449# a_1500_28546# 0.217f
C490 a_n1558_n8534# w_n1594_n8634# 0.0187f
C491 a_n1500_21033# a_1500_21130# 0.217f
C492 w_n1594_n60546# a_n1558_n60446# 0.0187f
C493 w_n1594_n28410# a_1500_n29546# 0.0023f
C494 w_n1594_n7398# a_n1500_n6159# 0.0172f
C495 w_n1594_n27174# a_n1558_n25838# 0.0023f
C496 a_n1558_47086# w_n1594_45750# 0.0023f
C497 w_n1594_27210# a_n1500_27213# 1.65f
C498 a_n1558_n49322# w_n1594_n48186# 0.0023f
C499 a_n1500_58113# a_n1500_56877# 3.11f
C500 w_n1594_29682# a_n1558_31018# 0.0023f
C501 a_1500_n33254# a_1500_n34490# 0.0105f
C502 a_n1558_32254# w_n1594_33390# 0.0023f
C503 a_1500_10006# w_n1594_8670# 0.0023f
C504 a_n1500_n34587# a_n1558_n34490# 0.217f
C505 w_n1594_42042# a_n1500_43281# 0.0172f
C506 a_n1500_n59307# a_1500_n59210# 0.217f
C507 w_n1594_n4926# a_n1558_n4826# 0.0187f
C508 a_n1500_n1215# a_1500_n1118# 0.217f
C509 a_n1558_58210# a_n1558_59446# 0.0105f
C510 a_n1558_n55502# a_n1558_n56738# 0.0105f
C511 w_n1594_13614# a_1500_14950# 0.0023f
C512 a_n1558_n17186# a_n1558_n18422# 0.0105f
C513 a_1500_12478# w_n1594_11142# 0.0023f
C514 w_n1594_38334# a_n1500_38337# 1.65f
C515 a_n1500_n27171# a_n1500_n28407# 3.11f
C516 a_n1500_51933# a_n1558_52030# 0.217f
C517 a_1500_53266# a_1500_52030# 0.0105f
C518 w_n1594_n32118# a_n1500_n32115# 1.65f
C519 a_n1500_60585# a_n1558_60682# 0.217f
C520 a_n1558_n54266# w_n1594_n53130# 0.0023f
C521 a_n1500_n50655# w_n1594_n51894# 0.0172f
C522 a_n1500_n43239# a_1500_n43142# 0.217f
C523 w_n1594_16086# a_n1558_16186# 0.0187f
C524 a_1500_n3590# w_n1594_n2454# 0.0023f
C525 w_n1594_n20994# a_1500_n22130# 0.0023f
C526 a_n1500_n20991# w_n1594_n19758# 0.0172f
C527 a_1500_8770# w_n1594_7434# 0.0023f
C528 w_n1594_48222# a_1500_47086# 0.0023f
C529 a_n1500_2493# a_n1558_2590# 0.217f
C530 a_n1558_18658# a_n1558_17422# 0.0105f
C531 w_n1594_39570# a_1500_39670# 0.0187f
C532 a_n1558_n35726# w_n1594_n34590# 0.0023f
C533 a_1500_n49322# a_1500_n50558# 0.0105f
C534 w_n1594_n58074# a_1500_n57974# 0.0187f
C535 a_n1500_n50655# a_n1558_n50558# 0.217f
C536 w_n1594_17322# a_n1500_16089# 0.0172f
C537 a_1500_n19658# a_1500_n20894# 0.0105f
C538 a_n1500_n12339# a_n1558_n12242# 0.217f
C539 a_1500_n11006# a_1500_n12242# 0.0105f
C540 w_n1594_n25938# a_n1558_n24602# 0.0023f
C541 a_n1558_45850# a_n1558_44614# 0.0105f
C542 w_n1594_1254# a_1500_118# 0.0023f
C543 a_1500_n46850# w_n1594_n45714# 0.0023f
C544 a_n1500_44517# w_n1594_43278# 0.0172f
C545 w_n1594_44514# a_n1500_43281# 0.0172f
C546 a_1500_n44378# w_n1594_n44478# 0.0187f
C547 w_n1594_n55602# a_1500_n55502# 0.0187f
C548 a_n1500_7437# w_n1594_6198# 0.0172f
C549 a_n1558_n3590# a_n1558_n4826# 0.0105f
C550 a_n1500_60585# w_n1594_59346# 0.0172f
C551 a_n1558_n40670# w_n1594_n39534# 0.0023f
C552 a_n1500_55641# w_n1594_55638# 1.65f
C553 a_n1500_3729# w_n1594_4962# 0.0172f
C554 a_n1558_55738# w_n1594_56874# 0.0023f
C555 a_n1500_n37059# w_n1594_n38298# 0.0172f
C556 a_n1500_8673# a_n1500_7437# 3.11f
C557 a_1500_32254# a_1500_31018# 0.0105f
C558 a_n1500_30921# a_n1558_31018# 0.217f
C559 a_n1500_23505# a_n1558_23602# 0.217f
C560 a_1500_24838# a_1500_23602# 0.0105f
C561 a_1500_n44378# a_1500_n45614# 0.0105f
C562 a_1500_n51794# w_n1594_n50658# 0.0023f
C563 w_n1594_n29646# a_n1558_n29546# 0.0187f
C564 a_n1558_n48086# w_n1594_n49422# 0.0023f
C565 w_n1594_n1218# a_n1558_n1118# 0.0187f
C566 w_n1594_46986# a_1500_48322# 0.0023f
C567 w_n1594_22266# a_n1558_23602# 0.0023f
C568 w_n1594_n23466# a_n1558_n22130# 0.0023f
C569 a_1500_33490# a_n1500_33393# 0.217f
C570 a_n1500_14853# a_1500_14950# 0.217f
C571 a_n1500_n13575# w_n1594_n14814# 0.0172f
C572 w_n1594_37098# a_n1500_35865# 0.0172f
C573 a_n1500_n9867# w_n1594_n11106# 0.0172f
C574 a_n1558_31018# w_n1594_32154# 0.0023f
C575 w_n1594_18# a_1500_1354# 0.0023f
C576 a_n1500_n24699# a_1500_n24602# 0.217f
C577 w_n1594_n6162# a_n1558_n7298# 0.0023f
C578 a_n1500_42045# a_1500_42142# 0.217f
C579 a_n1500_32157# w_n1594_30918# 0.0172f
C580 a_n1500_n40767# a_n1558_n40670# 0.217f
C581 w_n1594_35862# a_n1558_35962# 0.0187f
C582 a_1500_n39434# a_1500_n40670# 0.0105f
C583 w_n1594_49458# a_n1558_48322# 0.0023f
C584 a_n1500_n43239# w_n1594_n42006# 0.0172f
C585 a_n1500_35865# a_n1500_34629# 3.11f
C586 w_n1594_51930# a_n1558_52030# 0.0187f
C587 a_n1500_n7395# a_1500_n7298# 0.217f
C588 w_n1594_28446# a_n1500_29685# 0.0172f
C589 a_1500_n12242# w_n1594_n13578# 0.0023f
C590 a_n1500_58113# w_n1594_56874# 0.0172f
C591 a_1500_n38198# w_n1594_n37062# 0.0023f
C592 w_n1594_46986# a_n1500_48225# 0.0172f
C593 a_n1558_n34490# w_n1594_n35826# 0.0023f
C594 a_n1558_n17186# w_n1594_n18522# 0.0023f
C595 a_1500_59446# a_n1500_59349# 0.217f
C596 w_n1594_n60546# a_n1500_n61779# 0.0172f
C597 w_n1594_n7398# a_1500_n6062# 0.0023f
C598 w_n1594_n27174# a_n1500_n27171# 1.65f
C599 a_n1500_n14811# w_n1594_n16050# 0.0172f
C600 w_n1594_18558# a_n1500_19797# 0.0172f
C601 a_n1500_n45711# a_n1558_n45614# 0.217f
C602 a_n1500_45753# w_n1594_45750# 1.65f
C603 w_n1594_27210# a_1500_27310# 0.0187f
C604 a_1500_n45614# w_n1594_n46950# 0.0023f
C605 w_n1594_29682# a_n1500_29685# 1.65f
C606 w_n1594_42042# a_1500_43378# 0.0023f
C607 a_n1558_8770# w_n1594_8670# 0.0187f
C608 a_n1500_n34587# a_n1500_n35823# 3.11f
C609 w_n1594_n4926# a_n1500_n6159# 0.0172f
C610 w_n1594_23502# a_n1558_24838# 0.0023f
C611 a_n1500_n56835# a_n1558_n56738# 0.217f
C612 a_n1558_n19658# w_n1594_n20994# 0.0023f
C613 a_1500_n17186# a_1500_n18422# 0.0105f
C614 a_n1500_11145# a_1500_11242# 0.217f
C615 a_n1500_n18519# a_n1558_n18422# 0.217f
C616 a_n1558_11242# w_n1594_11142# 0.0187f
C617 w_n1594_38334# a_1500_38434# 0.0187f
C618 a_n1558_n27074# a_n1558_n28310# 0.0105f
C619 a_n1500_51933# a_n1500_50697# 3.11f
C620 w_n1594_n32118# a_1500_n32018# 0.0187f
C621 a_1500_n50558# w_n1594_n51894# 0.0023f
C622 a_n1558_58210# w_n1594_59346# 0.0023f
C623 w_n1594_16086# a_n1500_14853# 0.0172f
C624 a_1500_n33254# w_n1594_n32118# 0.0023f
C625 a_n1558_7534# w_n1594_7434# 0.0187f
C626 a_n1558_59446# w_n1594_60582# 0.0023f
C627 a_n1500_48225# a_1500_48322# 0.217f
C628 a_1500_18658# a_1500_17422# 0.0105f
C629 w_n1594_39570# a_n1558_38434# 0.0023f
C630 a_n1500_17325# a_n1558_17422# 0.217f
C631 a_n1500_n50655# a_n1500_n51891# 3.11f
C632 w_n1594_n58074# a_n1558_n59210# 0.0023f
C633 w_n1594_17322# a_1500_16186# 0.0023f
C634 a_n1500_n12339# a_n1500_n13575# 3.11f
C635 w_n1594_n25938# a_n1500_n25935# 1.65f
C636 a_n1500_44517# a_n1558_44614# 0.217f
C637 w_n1594_n22230# a_n1558_n22130# 0.0187f
C638 w_n1594_2490# a_1500_2590# 0.0187f
C639 a_1500_45850# a_1500_44614# 0.0105f
C640 a_n1500_n22227# a_n1558_n22130# 0.217f
C641 a_n1500_n56835# a_1500_n56738# 0.217f
C642 a_1500_44614# w_n1594_43278# 0.0023f
C643 w_n1594_44514# a_1500_43378# 0.0023f
C644 w_n1594_n55602# a_n1558_n56738# 0.0023f
C645 a_n1500_n42003# w_n1594_n43242# 0.0172f
C646 w_n1594_n54366# a_n1500_n53127# 0.0172f
C647 a_1500_13714# w_n1594_12378# 0.0023f
C648 a_n1500_38337# a_1500_38434# 0.217f
C649 a_1500_n3590# a_1500_n4826# 0.0105f
C650 a_1500_7534# w_n1594_6198# 0.0023f
C651 a_n1500_n4923# a_n1558_n4826# 0.217f
C652 a_1500_3826# w_n1594_4962# 0.0023f
C653 a_1500_n36962# w_n1594_n38298# 0.0023f
C654 a_1500_55738# w_n1594_55638# 0.0187f
C655 a_n1558_55738# w_n1594_54402# 0.0023f
C656 a_n1558_8770# a_n1558_7534# 0.0105f
C657 a_n1500_30921# a_n1500_29685# 3.11f
C658 w_n1594_n61782# a_n1500_n60543# 0.0172f
C659 a_n1500_n30879# a_1500_n30782# 0.217f
C660 a_n1500_23505# a_n1500_22269# 3.11f
C661 w_n1594_n29646# a_n1500_n30879# 0.0172f
C662 a_n1500_n49419# w_n1594_n49422# 1.65f
C663 a_n1500_55641# a_1500_55738# 0.217f
C664 w_n1594_n1218# a_n1500_n2451# 0.0172f
C665 w_n1594_46986# a_n1558_47086# 0.0187f
C666 w_n1594_n23466# a_n1500_n23463# 1.65f
C667 w_n1594_22266# a_n1500_22269# 1.65f
C668 a_1500_n13478# w_n1594_n14814# 0.0023f
C669 w_n1594_37098# a_1500_35962# 0.0023f
C670 a_1500_n9770# w_n1594_n11106# 0.0023f
C671 a_n1500_n16047# w_n1594_n17286# 0.0172f
C672 a_1500_39670# w_n1594_40806# 0.0023f
C673 w_n1594_n55602# a_1500_n56738# 0.0023f
C674 a_n1500_3729# w_n1594_2490# 0.0172f
C675 a_1500_32254# w_n1594_30918# 0.0023f
C676 a_n1558_5062# w_n1594_3726# 0.0023f
C677 a_n1500_21# a_1500_118# 0.217f
C678 w_n1594_35862# a_n1500_34629# 0.0172f
C679 w_n1594_34626# a_n1500_35865# 0.0172f
C680 a_n1500_n40767# a_n1500_n42003# 3.11f
C681 a_1500_n43142# w_n1594_n42006# 0.0023f
C682 a_n1558_35962# a_n1558_34726# 0.0105f
C683 w_n1594_51930# a_n1500_50697# 0.0172f
C684 w_n1594_28446# a_1500_29782# 0.0023f
C685 a_n1558_n39434# w_n1594_n40770# 0.0023f
C686 a_1500_40906# a_1500_39670# 0.0105f
C687 a_n1558_n13478# w_n1594_n13578# 0.0187f
C688 a_n1500_42045# w_n1594_40806# 0.0172f
C689 a_n1500_4965# a_1500_5062# 0.217f
C690 a_n1500_n35823# w_n1594_n35826# 1.65f
C691 a_n1500_n18519# w_n1594_n18522# 1.65f
C692 a_n1500_n9867# a_n1500_n8631# 3.11f
C693 w_n1594_n60546# a_1500_n61682# 0.0023f
C694 w_n1594_9906# a_n1500_11145# 0.0172f
C695 w_n1594_n59310# a_n1558_n57974# 0.0023f
C696 w_n1594_n7398# a_n1558_n7298# 0.0187f
C697 w_n1594_n27174# a_1500_n27074# 0.0187f
C698 a_n1500_n48183# a_1500_n48086# 0.217f
C699 a_n1500_n9867# a_1500_n9770# 0.217f
C700 w_n1594_18558# a_1500_19894# 0.0023f
C701 a_1500_n14714# w_n1594_n16050# 0.0023f
C702 a_n1500_n45711# a_n1500_n46947# 3.11f
C703 a_1500_45850# w_n1594_45750# 0.0187f
C704 w_n1594_27210# a_n1558_26074# 0.0023f
C705 a_n1558_n46850# w_n1594_n46950# 0.0187f
C706 a_n1558_n44378# w_n1594_n45714# 0.0023f
C707 a_n1558_n34490# a_n1558_n35726# 0.0105f
C708 w_n1594_29682# a_1500_29782# 0.0187f
C709 w_n1594_42042# a_n1558_42142# 0.0187f
C710 a_n1500_7437# w_n1594_8670# 0.0172f
C711 w_n1594_n56838# a_n1558_n55502# 0.0023f
C712 w_n1594_n4926# a_1500_n6062# 0.0023f
C713 a_n1558_60682# w_n1594_60582# 0.0187f
C714 w_n1594_23502# a_n1500_23505# 1.65f
C715 a_n1500_n20991# w_n1594_n20994# 1.65f
C716 a_n1500_n18519# a_n1500_n19755# 3.11f
C717 w_n1594_38334# a_n1558_37198# 0.0023f
C718 a_n1500_9909# w_n1594_11142# 0.0172f
C719 a_n1500_n28407# a_n1558_n28310# 0.217f
C720 a_1500_n27074# a_1500_n28310# 0.0105f
C721 a_n1558_52030# a_n1558_50794# 0.0105f
C722 a_n1558_n51794# w_n1594_n51894# 0.0187f
C723 w_n1594_n30882# a_n1500_n29643# 0.0172f
C724 w_n1594_16086# a_1500_14950# 0.0023f
C725 a_n1500_34629# w_n1594_33390# 0.0172f
C726 w_n1594_n33354# a_n1558_n32018# 0.0023f
C727 a_n1558_59446# w_n1594_58110# 0.0023f
C728 a_n1500_6201# w_n1594_7434# 0.0172f
C729 a_n1500_17325# a_n1500_16089# 3.11f
C730 a_n1558_n33254# w_n1594_n33354# 0.0187f
C731 a_n1558_n50558# a_n1558_n51794# 0.0105f
C732 w_n1594_21030# a_n1558_22366# 0.0023f
C733 a_n1558_n12242# a_n1558_n13478# 0.0105f
C734 w_n1594_n25938# a_1500_n25838# 0.0187f
C735 a_n1500_n22227# a_n1500_n23463# 3.11f
C736 a_n1500_44517# a_n1500_43281# 3.11f
C737 w_n1594_3726# a_1500_2590# 0.0023f
C738 w_n1594_2490# a_n1558_1354# 0.0023f
C739 w_n1594_n22230# a_n1500_n23463# 0.0172f
C740 a_n1558_43378# w_n1594_43278# 0.0187f
C741 a_n1500_n38295# a_1500_n38198# 0.217f
C742 a_1500_n41906# w_n1594_n43242# 0.0023f
C743 w_n1594_n54366# a_1500_n53030# 0.0023f
C744 w_n1594_39570# a_n1558_40906# 0.0023f
C745 a_n1558_12478# w_n1594_12378# 0.0187f
C746 a_n1558_6298# w_n1594_6198# 0.0187f
C747 a_n1500_n4923# a_n1500_n6159# 3.11f
C748 a_n1558_n38198# w_n1594_n38298# 0.0187f
C749 a_n1558_54502# w_n1594_55638# 0.0023f
C750 a_n1500_54405# w_n1594_54402# 1.65f
C751 a_1500_8770# a_1500_7534# 0.0105f
C752 a_n1500_7437# a_n1558_7534# 0.217f
C753 a_n1558_31018# a_n1558_29782# 0.0105f
C754 w_n1594_n61782# a_1500_n60446# 0.0023f
C755 a_n1558_23602# a_n1558_22366# 0.0105f
C756 a_n1500_53169# w_n1594_54402# 0.0172f
C757 a_1500_n49322# w_n1594_n49422# 0.0187f
C758 w_n1594_n29646# a_1500_n30782# 0.0023f
C759 w_n1594_n1218# a_1500_n2354# 0.0023f
C760 a_n1558_58210# a_n1558_56974# 0.0105f
C761 w_n1594_46986# a_n1500_45753# 0.0172f
C762 w_n1594_n23466# a_1500_n23366# 0.0187f
C763 w_n1594_22266# a_1500_22366# 0.0187f
C764 a_n1558_n14714# w_n1594_n14814# 0.0187f
C765 w_n1594_39570# a_1500_40906# 0.0023f
C766 a_n1558_n11006# w_n1594_n11106# 0.0187f
C767 a_n1500_n54363# a_1500_n54266# 0.217f
C768 a_1500_n15950# w_n1594_n17286# 0.0023f
C769 a_n1500_n16047# a_1500_n15950# 0.217f
C770 w_n1594_n3690# a_n1500_n2451# 0.0172f
C771 a_1500_3826# w_n1594_2490# 0.0023f
C772 a_n1500_3729# w_n1594_3726# 1.65f
C773 a_n1558_31018# w_n1594_30918# 0.0187f
C774 a_n1558_n40670# a_n1558_n41906# 0.0105f
C775 w_n1594_34626# a_1500_35962# 0.0023f
C776 w_n1594_35862# a_1500_34726# 0.0023f
C777 a_1500_35962# a_1500_34726# 0.0105f
C778 a_n1500_34629# a_n1558_34726# 0.217f
C779 a_n1500_n40767# w_n1594_n40770# 1.65f
C780 w_n1594_51930# a_1500_50794# 0.0023f
C781 w_n1594_28446# a_n1558_28546# 0.0187f
C782 a_n1500_n14811# w_n1594_n13578# 0.0172f
C783 a_1500_42142# w_n1594_40806# 0.0023f
C784 a_n1500_27213# a_1500_27310# 0.217f
C785 a_n1500_19797# a_1500_19894# 0.217f
C786 a_1500_n18422# w_n1594_n18522# 0.0187f
C787 a_1500_n35726# w_n1594_n35826# 0.0187f
C788 a_n1500_33393# w_n1594_32154# 0.0172f
C789 a_n1558_n9770# a_n1558_n8534# 0.0105f
C790 w_n1594_9906# a_1500_11242# 0.0023f
C791 w_n1594_25974# a_n1558_27310# 0.0023f
C792 w_n1594_n27174# a_n1558_n28310# 0.0023f
C793 w_n1594_n7398# a_n1500_n8631# 0.0172f
C794 w_n1594_n59310# a_n1500_n59307# 1.65f
C795 w_n1594_18558# a_n1558_18658# 0.0187f
C796 a_n1558_n15950# w_n1594_n16050# 0.0187f
C797 a_n1558_44614# w_n1594_45750# 0.0023f
C798 a_n1500_46989# a_1500_47086# 0.217f
C799 a_n1500_n48183# w_n1594_n46950# 0.0172f
C800 a_1500_42142# a_1500_40906# 0.0105f
C801 a_n1500_n35823# a_n1558_n35726# 0.217f
C802 a_1500_n34490# a_1500_n35726# 0.0105f
C803 w_n1594_29682# a_n1558_28546# 0.0023f
C804 a_1500_7534# w_n1594_8670# 0.0023f
C805 w_n1594_42042# a_n1500_40809# 0.0172f
C806 w_n1594_n56838# a_n1500_n56835# 1.65f
C807 w_n1594_18# a_1500_118# 0.0187f
C808 a_n1500_n60543# a_1500_n60446# 0.217f
C809 w_n1594_23502# a_1500_23602# 0.0187f
C810 a_n1500_n2451# a_1500_n2354# 0.217f
C811 a_n1500_21# a_n1500_n1215# 3.11f
C812 a_n1558_n18422# a_n1558_n19658# 0.0105f
C813 a_1500_10006# w_n1594_11142# 0.0023f
C814 a_n1500_n28407# a_n1500_n29643# 3.11f
C815 a_n1500_50697# a_n1558_50794# 0.217f
C816 a_1500_52030# a_1500_50794# 0.0105f
C817 a_n1558_n9770# w_n1594_n9870# 0.0187f
C818 a_n1500_n11103# w_n1594_n12342# 0.0172f
C819 a_n1500_n44475# a_1500_n44378# 0.217f
C820 w_n1594_n30882# a_1500_n29546# 0.0023f
C821 a_n1500_n53127# w_n1594_n51894# 0.0172f
C822 a_1500_34726# w_n1594_33390# 0.0023f
C823 w_n1594_n33354# a_n1500_n33351# 1.65f
C824 w_n1594_19794# a_n1558_21130# 0.0023f
C825 a_1500_6298# w_n1594_7434# 0.0023f
C826 a_n1558_17422# a_n1558_16186# 0.0105f
C827 a_n1500_n34587# w_n1594_n33354# 0.0172f
C828 a_1500_n50558# a_1500_n51794# 0.0105f
C829 a_n1500_n51891# a_n1558_n51794# 0.217f
C830 a_1500_n12242# a_1500_n13478# 0.0105f
C831 a_n1500_n13575# a_n1558_n13478# 0.217f
C832 w_n1594_21030# a_n1500_21033# 1.65f
C833 w_n1594_n25938# a_n1558_n27074# 0.0023f
C834 a_n1558_44614# a_n1558_43378# 0.0105f
C835 w_n1594_n22230# a_1500_n23366# 0.0023f
C836 w_n1594_n24702# a_n1500_n23463# 0.0172f
C837 a_n1558_n22130# a_n1558_n23366# 0.0105f
C838 a_n1558_n45614# w_n1594_n44478# 0.0023f
C839 a_n1500_42045# w_n1594_43278# 0.0172f
C840 a_n1500_n45711# w_n1594_n45714# 1.65f
C841 a_n1558_n43142# w_n1594_n43242# 0.0187f
C842 a_n1500_11145# w_n1594_12378# 0.0172f
C843 w_n1594_50694# a_n1558_52030# 0.0023f
C844 w_n1594_n54366# a_n1558_n54266# 0.0187f
C845 a_n1558_n4826# a_n1558_n6062# 0.0105f
C846 a_n1500_4965# w_n1594_6198# 0.0172f
C847 a_n1500_39573# a_n1558_39670# 0.217f
C848 a_n1500_n39531# w_n1594_n38298# 0.0172f
C849 a_1500_54502# w_n1594_54402# 0.0187f
C850 a_n1500_29685# a_n1558_29782# 0.217f
C851 a_1500_31018# a_1500_29782# 0.0105f
C852 a_n1500_7437# a_n1500_6201# 3.11f
C853 w_n1594_14850# a_1500_13714# 0.0023f
C854 a_n1500_22269# a_n1558_22366# 0.217f
C855 w_n1594_n61782# a_n1558_n61682# 0.0187f
C856 a_1500_23602# a_1500_22366# 0.0105f
C857 a_n1500_24741# a_1500_24838# 0.217f
C858 w_n1594_n28410# a_n1558_n27074# 0.0023f
C859 a_1500_53266# w_n1594_54402# 0.0023f
C860 a_1500_59446# w_n1594_60582# 0.0023f
C861 a_n1558_n50558# w_n1594_n49422# 0.0023f
C862 a_n1500_n46947# w_n1594_n48186# 0.0172f
C863 w_n1594_46986# a_1500_45850# 0.0023f
C864 w_n1594_22266# a_n1558_21130# 0.0023f
C865 w_n1594_n23466# a_n1558_n24602# 0.0023f
C866 a_n1500_n58071# a_n1558_n57974# 0.217f
C867 a_1500_n56738# a_1500_n57974# 0.0105f
C868 a_n1500_n16047# w_n1594_n14814# 0.0172f
C869 w_n1594_1254# a_1500_2590# 0.0023f
C870 a_n1500_54405# a_n1500_53169# 3.11f
C871 a_n1500_n12339# w_n1594_n11106# 0.0172f
C872 a_n1558_n17186# w_n1594_n17286# 0.0187f
C873 w_n1594_n3690# a_1500_n2354# 0.0023f
C874 a_n1558_13714# a_n1558_12478# 0.0105f
C875 a_n1500_n25935# a_1500_n25838# 0.217f
C876 w_n1594_14850# a_n1500_16089# 0.0172f
C877 a_n1500_29685# w_n1594_30918# 0.0172f
C878 a_n1558_2590# w_n1594_2490# 0.0187f
C879 a_1500_3826# w_n1594_3726# 0.0187f
C880 a_1500_58210# w_n1594_58110# 0.0187f
C881 a_n1500_n51891# w_n1594_n53130# 0.0172f
C882 a_n1500_n42003# a_n1558_n41906# 0.217f
C883 a_1500_n40670# a_1500_n41906# 0.0105f
C884 w_n1594_34626# a_n1558_34726# 0.0187f
C885 a_n1558_n1118# w_n1594_n2454# 0.0023f
C886 a_n1500_34629# a_n1500_33393# 3.11f
C887 w_n1594_28446# a_n1500_27213# 0.0172f
C888 a_n1500_n8631# a_1500_n8534# 0.217f
C889 a_1500_n40670# w_n1594_n40770# 0.0187f
C890 a_1500_n14714# w_n1594_n13578# 0.0023f
C891 a_n1558_40906# w_n1594_40806# 0.0187f
C892 a_n1558_n19658# w_n1594_n18522# 0.0023f
C893 a_1500_n9770# a_1500_n8534# 0.0105f
C894 a_n1558_n36962# w_n1594_n35826# 0.0023f
C895 w_n1594_n59310# a_1500_n59210# 0.0187f
C896 w_n1594_9906# a_n1558_10006# 0.0187f
C897 w_n1594_n7398# a_1500_n8534# 0.0023f
C898 w_n1594_25974# a_n1500_25977# 1.65f
C899 w_n1594_18558# a_n1500_17325# 0.0172f
C900 a_n1500_n17283# w_n1594_n16050# 0.0172f
C901 a_1500_n48086# w_n1594_n46950# 0.0023f
C902 a_n1500_n35823# a_n1500_n37059# 3.11f
C903 w_n1594_25974# a_n1558_24838# 0.0023f
C904 w_n1594_23502# a_n1558_22366# 0.0023f
C905 a_n1500_n38295# w_n1594_n39534# 0.0172f
C906 a_1500_n18422# a_1500_n19658# 0.0105f
C907 a_n1500_n19755# a_n1558_n19658# 0.217f
C908 w_n1594_n9870# a_n1558_n8534# 0.0023f
C909 a_n1500_9909# a_1500_10006# 0.217f
C910 w_n1594_38334# a_n1500_39573# 0.0172f
C911 a_1500_40906# w_n1594_40806# 0.0187f
C912 a_n1558_n28310# a_n1558_n29546# 0.0105f
C913 a_n1500_50697# a_n1500_49461# 3.11f
C914 a_1500_n11006# w_n1594_n12342# 0.0023f
C915 a_n1500_n11103# w_n1594_n9870# 0.0172f
C916 w_n1594_n30882# a_n1558_n30782# 0.0187f
C917 a_1500_n53030# w_n1594_n51894# 0.0023f
C918 a_n1558_n49322# w_n1594_n50658# 0.0023f
C919 a_n1558_33490# w_n1594_33390# 0.0187f
C920 a_n1558_n20894# w_n1594_n22230# 0.0023f
C921 w_n1594_19794# a_n1500_19797# 1.65f
C922 a_1500_17422# a_1500_16186# 0.0105f
C923 a_n1500_16089# a_n1558_16186# 0.217f
C924 a_1500_n34490# w_n1594_n33354# 0.0023f
C925 a_n1500_n51891# a_n1500_n53127# 3.11f
C926 a_n1500_n13575# a_n1500_n14811# 3.11f
C927 w_n1594_n56838# a_n1500_n58071# 0.0172f
C928 w_n1594_24738# a_n1500_25977# 0.0172f
C929 w_n1594_21030# a_1500_21130# 0.0187f
C930 w_n1594_18# a_n1500_n1215# 0.0172f
C931 w_n1594_n6162# a_n1500_n4923# 0.0172f
C932 a_n1500_60585# a_n1500_59349# 3.11f
C933 a_n1500_n23463# a_n1558_n23366# 0.217f
C934 a_1500_n22130# a_1500_n23366# 0.0105f
C935 a_n1500_43281# a_n1558_43378# 0.217f
C936 w_n1594_n24702# a_1500_n23366# 0.0023f
C937 a_1500_44614# a_1500_43378# 0.0105f
C938 a_1500_42142# w_n1594_43278# 0.0023f
C939 a_n1500_n44475# w_n1594_n43242# 0.0172f
C940 w_n1594_49458# a_n1500_50697# 0.0172f
C941 a_1500_13714# w_n1594_13614# 0.0187f
C942 a_n1500_37101# a_1500_37198# 0.217f
C943 w_n1594_n54366# a_n1500_n55599# 0.0172f
C944 a_1500_n4826# a_1500_n6062# 0.0105f
C945 a_1500_11242# w_n1594_12378# 0.0023f
C946 w_n1594_50694# a_n1500_50697# 1.65f
C947 a_n1500_n6159# a_n1558_n6062# 0.217f
C948 a_1500_5062# w_n1594_6198# 0.0023f
C949 a_n1500_39573# a_n1500_38337# 3.11f
C950 a_1500_n39434# w_n1594_n38298# 0.0023f
C951 w_n1594_24738# a_n1558_24838# 0.0187f
C952 a_1500_3826# a_1500_2590# 0.0105f
C953 a_n1500_29685# a_n1500_28449# 3.11f
C954 a_n1558_7534# a_n1558_6298# 0.0105f
C955 a_n1558_n35726# w_n1594_n37062# 0.0023f
C956 a_n1500_n32115# a_1500_n32018# 0.217f
C957 a_n1500_22269# a_n1500_21033# 3.11f
C958 w_n1594_n28410# a_n1500_n28407# 1.65f
C959 a_n1558_n45614# a_n1558_n46850# 0.0105f
C960 a_n1558_n33254# a_n1558_n32018# 0.0105f
C961 a_1500_59446# w_n1594_58110# 0.0023f
C962 a_n1500_54405# a_1500_54502# 0.217f
C963 a_1500_n46850# w_n1594_n48186# 0.0023f
C964 a_1500_n15950# w_n1594_n14814# 0.0023f
C965 a_1500_60682# w_n1594_59346# 0.0023f
C966 a_n1558_54502# a_n1558_53266# 0.0105f
C967 a_1500_n12242# w_n1594_n11106# 0.0023f
C968 a_n1500_n58071# a_n1500_n59307# 3.11f
C969 w_n1594_1254# a_n1558_1354# 0.0187f
C970 a_n1500_n18519# w_n1594_n17286# 0.0172f
C971 a_1500_13714# a_1500_12478# 0.0105f
C972 w_n1594_12378# a_n1500_13617# 0.0172f
C973 w_n1594_n3690# a_n1558_n3590# 0.0187f
C974 a_n1500_12381# a_n1558_12478# 0.217f
C975 a_1500_29782# w_n1594_30918# 0.0023f
C976 w_n1594_14850# a_1500_16186# 0.0023f
C977 a_n1500_53169# a_1500_53266# 0.217f
C978 a_n1558_2590# w_n1594_3726# 0.0023f
C979 a_1500_n51794# w_n1594_n53130# 0.0023f
C980 a_n1558_56974# w_n1594_58110# 0.0023f
C981 a_n1500_n42003# a_n1500_n43239# 3.11f
C982 w_n1594_34626# a_n1500_33393# 0.0172f
C983 a_n1558_34726# a_n1558_33490# 0.0105f
C984 a_n1500_n2451# w_n1594_n2454# 1.65f
C985 w_n1594_28446# a_1500_27310# 0.0023f
C986 a_n1558_n41906# w_n1594_n40770# 0.0023f
C987 a_n1558_n18422# w_n1594_n19758# 0.0023f
C988 a_n1500_3729# a_1500_3826# 0.217f
C989 a_1500_n33254# w_n1594_n34590# 0.0023f
C990 w_n1594_9906# a_n1500_8673# 0.0172f
C991 w_n1594_n59310# a_n1558_n60446# 0.0023f
C992 w_n1594_25974# a_1500_26074# 0.0187f
C993 a_n1500_n49419# a_1500_n49322# 0.217f
C994 w_n1594_18558# a_1500_17422# 0.0023f
C995 w_n1594_17322# a_n1558_18658# 0.0023f
C996 a_1500_n17186# w_n1594_n16050# 0.0023f
C997 a_n1500_n11103# a_1500_n11006# 0.217f
C998 a_n1558_13714# a_n1558_14950# 0.0105f
C999 w_n1594_44514# a_n1558_45850# 0.0023f
C1000 a_n1558_n35726# a_n1558_n36962# 0.0105f
C1001 a_n1500_n43239# w_n1594_n44478# 0.0172f
C1002 w_n1594_n55602# a_n1500_n54363# 0.0172f
C1003 a_n1558_6298# w_n1594_4962# 0.0023f
C1004 a_1500_n38198# w_n1594_n39534# 0.0023f
C1005 a_1500_58210# w_n1594_56874# 0.0023f
C1006 w_n1594_n22230# a_1500_n20894# 0.0023f
C1007 a_n1500_1257# a_1500_1354# 0.217f
C1008 a_n1500_n19755# a_n1500_n20991# 3.11f
C1009 a_n1500_32157# a_1500_32254# 0.217f
C1010 w_n1594_48222# a_n1558_49558# 0.0023f
C1011 a_1500_n28310# a_1500_n29546# 0.0105f
C1012 a_n1500_n29643# a_n1558_n29546# 0.217f
C1013 a_n1558_50794# a_n1558_49558# 0.0105f
C1014 a_1500_n11006# w_n1594_n9870# 0.0023f
C1015 a_n1558_n12242# w_n1594_n12342# 0.0187f
C1016 w_n1594_n30882# a_n1500_n32115# 0.0172f
C1017 a_n1500_n50655# w_n1594_n50658# 1.65f
C1018 a_1500_58210# a_1500_56974# 0.0105f
C1019 a_n1500_56877# a_n1558_56974# 0.217f
C1020 w_n1594_19794# a_1500_19894# 0.0187f
C1021 a_n1500_16089# a_n1500_14853# 3.11f
C1022 w_n1594_37098# a_n1558_38434# 0.0023f
C1023 a_n1558_54502# w_n1594_53166# 0.0023f
C1024 a_n1558_n51794# a_n1558_n53030# 0.0105f
C1025 w_n1594_n56838# a_1500_n57974# 0.0023f
C1026 w_n1594_24738# a_1500_26074# 0.0023f
C1027 a_n1558_n13478# a_n1558_n14714# 0.0105f
C1028 w_n1594_21030# a_n1558_19894# 0.0023f
C1029 w_n1594_18# a_1500_n1118# 0.0023f
C1030 w_n1594_n6162# a_1500_n4826# 0.0023f
C1031 a_n1500_n23463# a_n1500_n24699# 3.11f
C1032 a_1500_33490# w_n1594_32154# 0.0023f
C1033 a_n1500_43281# a_n1500_42045# 3.11f
C1034 w_n1594_n24702# a_n1558_n24602# 0.0187f
C1035 a_n1558_53266# w_n1594_53166# 0.0187f
C1036 a_n1500_n39531# a_1500_n39434# 0.217f
C1037 a_1500_n44378# w_n1594_n43242# 0.0023f
C1038 a_n1558_n40670# w_n1594_n42006# 0.0023f
C1039 w_n1594_49458# a_1500_50794# 0.0023f
C1040 a_n1500_n6159# a_n1500_n7395# 3.11f
C1041 w_n1594_50694# a_1500_50794# 0.0187f
C1042 a_n1558_12478# w_n1594_13614# 0.0023f
C1043 w_n1594_n54366# a_1500_n55502# 0.0023f
C1044 w_n1594_24738# a_n1500_23505# 0.0172f
C1045 a_n1500_6201# a_n1558_6298# 0.217f
C1046 a_1500_7534# a_1500_6298# 0.0105f
C1047 a_n1500_2493# a_n1500_1257# 3.11f
C1048 a_n1500_n37059# w_n1594_n37062# 1.65f
C1049 a_n1558_29782# a_n1558_28546# 0.0105f
C1050 a_n1558_n7298# w_n1594_n8634# 0.0023f
C1051 a_n1558_22366# a_n1558_21130# 0.0105f
C1052 w_n1594_n60546# a_n1558_n59210# 0.0023f
C1053 w_n1594_n28410# a_1500_n28310# 0.0187f
C1054 a_n1500_n46947# a_n1558_n46850# 0.217f
C1055 a_1500_n45614# a_1500_n46850# 0.0105f
C1056 a_n1500_n9867# w_n1594_n8634# 0.0172f
C1057 a_n1558_n33254# a_n1500_n33351# 0.217f
C1058 a_1500_n33254# a_1500_n32018# 0.0105f
C1059 w_n1594_27210# a_n1500_28449# 0.0172f
C1060 a_n1558_n48086# w_n1594_n48186# 0.0187f
C1061 a_n1500_40809# a_n1500_39573# 3.11f
C1062 w_n1594_n58074# a_n1558_n56738# 0.0023f
C1063 w_n1594_n4926# a_n1558_n3590# 0.0023f
C1064 w_n1594_1254# a_n1500_21# 0.0172f
C1065 a_1500_54502# a_1500_53266# 0.0105f
C1066 a_n1558_n57974# a_n1558_n59210# 0.0105f
C1067 a_n1500_n55599# a_1500_n55502# 0.217f
C1068 a_1500_n18422# w_n1594_n17286# 0.0023f
C1069 a_n1500_12381# a_n1500_11145# 3.11f
C1070 a_n1500_n17283# a_1500_n17186# 0.217f
C1071 w_n1594_n3690# a_n1500_n4923# 0.0172f
C1072 w_n1594_14850# a_n1558_14950# 0.0187f
C1073 w_n1594_n32118# a_n1500_n30879# 0.0172f
C1074 a_n1558_n53030# w_n1594_n53130# 0.0187f
C1075 a_n1558_n41906# a_n1558_n43142# 0.0105f
C1076 w_n1594_16086# a_n1558_17422# 0.0023f
C1077 a_1500_n2354# w_n1594_n2454# 0.0187f
C1078 a_n1500_33393# a_n1558_33490# 0.217f
C1079 a_n1500_n19755# w_n1594_n19758# 1.65f
C1080 a_n1500_25977# a_1500_26074# 0.217f
C1081 w_n1594_48222# a_1500_48322# 0.0187f
C1082 a_n1500_18561# a_1500_18658# 0.217f
C1083 a_n1558_n34490# w_n1594_n34590# 0.0187f
C1084 a_1500_59446# a_1500_60682# 0.0105f
C1085 w_n1594_n1218# a_1500_118# 0.0023f
C1086 w_n1594_9906# a_1500_8770# 0.0023f
C1087 w_n1594_n58074# a_1500_n56738# 0.0023f
C1088 w_n1594_17322# a_n1500_17325# 1.65f
C1089 a_1500_13714# a_1500_14950# 0.0105f
C1090 a_n1558_13714# a_n1500_13617# 0.217f
C1091 a_n1500_45753# a_1500_45850# 0.217f
C1092 a_1500_n45614# w_n1594_n45714# 0.0187f
C1093 w_n1594_44514# a_n1500_44517# 1.65f
C1094 a_n1500_n37059# a_n1558_n36962# 0.217f
C1095 a_1500_n43142# w_n1594_n44478# 0.0023f
C1096 a_1500_n35726# a_1500_n36962# 0.0105f
C1097 w_n1594_n55602# a_1500_n54266# 0.0023f
C1098 a_n1500_n61779# a_1500_n61682# 0.217f
C1099 a_n1500_n3687# a_1500_n3590# 0.217f
C1100 a_n1558_2590# w_n1594_1254# 0.0023f
C1101 w_n1594_23502# a_n1500_24741# 0.0172f
C1102 a_n1558_56974# w_n1594_56874# 0.0187f
C1103 a_1500_n20894# a_1500_n22130# 0.0105f
C1104 a_n1500_4965# w_n1594_4962# 1.65f
C1105 a_n1500_56877# w_n1594_55638# 0.0172f
C1106 a_n1558_n39434# w_n1594_n39534# 0.0187f
C1107 a_n1558_n19658# a_n1558_n20894# 0.0105f
C1108 a_n1500_n29643# a_n1500_n30879# 3.11f
C1109 w_n1594_48222# a_n1500_48225# 1.65f
C1110 a_1500_50794# a_1500_49558# 0.0105f
C1111 a_n1500_49461# a_n1558_49558# 0.217f
C1112 a_n1500_n13575# w_n1594_n12342# 0.0172f
C1113 w_n1594_n30882# a_1500_n32018# 0.0023f
C1114 w_n1594_n29646# a_n1558_n28310# 0.0023f
C1115 a_1500_n50558# w_n1594_n50658# 0.0187f
C1116 a_n1500_58113# w_n1594_59346# 0.0172f
C1117 a_n1500_56877# a_n1500_55641# 3.11f
C1118 w_n1594_19794# a_n1558_18658# 0.0023f
C1119 a_n1500_59349# w_n1594_60582# 0.0172f
C1120 a_n1558_16186# a_n1558_14950# 0.0105f
C1121 w_n1594_37098# a_n1500_37101# 1.65f
C1122 a_n1500_n53127# a_n1558_n53030# 0.217f
C1123 a_1500_n51794# a_1500_n53030# 0.0105f
C1124 a_n1500_n14811# a_n1558_n14714# 0.217f
C1125 a_1500_n13478# a_1500_n14714# 0.0105f
C1126 w_n1594_n6162# a_n1558_n6062# 0.0187f
C1127 w_n1594_n24702# a_n1500_n25935# 0.0172f
C1128 a_n1558_32254# w_n1594_32154# 0.0187f
C1129 a_n1558_n23366# a_n1558_n24602# 0.0105f
C1130 a_n1500_51933# w_n1594_53166# 0.0172f
C1131 a_n1558_43378# a_n1558_42142# 0.0105f
C1132 w_n1594_35862# a_n1558_37198# 0.0023f
C1133 w_n1594_49458# a_n1558_49558# 0.0187f
C1134 a_n1500_n42003# w_n1594_n42006# 1.65f
C1135 a_n1558_n6062# a_n1558_n7298# 0.0105f
C1136 w_n1594_50694# a_n1558_49558# 0.0023f
C1137 w_n1594_51930# a_n1558_53266# 0.0023f
C1138 w_n1594_24738# a_1500_23602# 0.0023f
C1139 a_1500_n36962# w_n1594_n37062# 0.0187f
C1140 a_1500_29782# a_1500_28546# 0.0105f
C1141 a_n1500_6201# a_n1500_4965# 3.11f
C1142 a_n1558_2590# a_n1558_1354# 0.0105f
C1143 a_n1500_28449# a_n1558_28546# 0.217f
C1144 a_n1500_n8631# w_n1594_n8634# 1.65f
C1145 a_1500_22366# a_1500_21130# 0.0105f
C1146 a_n1500_21033# a_n1558_21130# 0.217f
C1147 w_n1594_n60546# a_n1500_n60543# 1.65f
C1148 w_n1594_n28410# a_n1558_n29546# 0.0023f
C1149 a_n1500_n46947# a_n1500_n48183# 3.11f
C1150 w_n1594_n27174# a_n1500_n25935# 0.0172f
C1151 a_1500_n9770# w_n1594_n8634# 0.0023f
C1152 a_n1500_n34587# a_n1500_n33351# 3.11f
C1153 a_n1500_46989# w_n1594_45750# 0.0172f
C1154 a_n1500_n49419# w_n1594_n48186# 0.0172f
C1155 w_n1594_27210# a_1500_28546# 0.0023f
C1156 a_n1500_58113# a_1500_58210# 0.217f
C1157 w_n1594_29682# a_n1500_30921# 0.0172f
C1158 a_n1500_32157# w_n1594_33390# 0.0172f
C1159 a_n1558_10006# w_n1594_8670# 0.0023f
C1160 a_n1500_n59307# a_n1558_n59210# 0.217f
C1161 a_1500_n57974# a_1500_n59210# 0.0105f
C1162 w_n1594_n4926# a_n1500_n4923# 1.65f
C1163 a_n1500_n1215# a_n1558_n1118# 0.217f
C1164 w_n1594_n3690# a_1500_n4826# 0.0023f
C1165 w_n1594_13614# a_n1558_14950# 0.0023f
C1166 a_n1558_12478# a_n1558_11242# 0.0105f
C1167 a_n1558_12478# w_n1594_11142# 0.0023f
C1168 w_n1594_38334# a_1500_39670# 0.0023f
C1169 a_n1500_n27171# a_1500_n27074# 0.217f
C1170 w_n1594_14850# a_n1500_13617# 0.0172f
C1171 a_n1500_n54363# w_n1594_n53130# 0.0172f
C1172 w_n1594_n32118# a_1500_n30782# 0.0023f
C1173 a_n1500_n43239# a_n1558_n43142# 0.217f
C1174 a_1500_n41906# a_1500_n43142# 0.0105f
C1175 w_n1594_16086# a_n1500_16089# 1.65f
C1176 a_n1558_n3590# w_n1594_n2454# 0.0023f
C1177 w_n1594_n20994# a_n1558_n22130# 0.0023f
C1178 a_1500_n19658# w_n1594_n19758# 0.0187f
C1179 w_n1594_48222# a_n1558_47086# 0.0023f
C1180 a_n1558_8770# w_n1594_7434# 0.0023f
C1181 w_n1594_39570# a_n1558_39670# 0.0187f
C1182 a_n1500_n35823# w_n1594_n34590# 0.0172f
C1183 w_n1594_n58074# a_n1558_n57974# 0.0187f
C1184 w_n1594_17322# a_1500_17422# 0.0187f
C1185 w_n1594_n25938# a_n1500_n24699# 0.0172f
C1186 w_n1594_1254# a_n1558_118# 0.0023f
C1187 a_n1500_12381# a_n1500_13617# 3.11f
C1188 a_n1558_n46850# w_n1594_n45714# 0.0023f
C1189 w_n1594_44514# a_1500_44614# 0.0187f
C1190 a_n1500_n37059# a_n1500_n38295# 3.11f
C1191 a_n1558_n44378# w_n1594_n44478# 0.0187f
C1192 w_n1594_n55602# a_n1558_n55502# 0.0187f
C1193 a_n1558_39670# a_n1558_38434# 0.0105f
C1194 a_n1500_60585# w_n1594_60582# 1.65f
C1195 a_n1500_n40767# w_n1594_n39534# 0.0172f
C1196 a_n1500_55641# w_n1594_56874# 0.0172f
C1197 a_1500_5062# w_n1594_4962# 0.0187f
C1198 a_1500_56974# w_n1594_55638# 0.0023f
C1199 a_n1500_8673# a_1500_8770# 0.217f
C1200 a_n1500_n20991# a_n1558_n20894# 0.217f
C1201 a_n1558_n29546# a_n1558_n30782# 0.0105f
C1202 a_n1500_49461# a_n1500_48225# 3.11f
C1203 a_1500_n13478# w_n1594_n12342# 0.0023f
C1204 w_n1594_49458# a_1500_48322# 0.0023f
C1205 a_n1558_n51794# w_n1594_n50658# 0.0023f
C1206 w_n1594_n29646# a_n1500_n29643# 1.65f
C1207 a_n1500_n48183# w_n1594_n49422# 0.0172f
C1208 w_n1594_n1218# a_n1500_n1215# 1.65f
C1209 a_n1558_56974# a_n1558_55738# 0.0105f
C1210 w_n1594_22266# a_n1500_23505# 0.0172f
C1211 w_n1594_n23466# a_n1500_n22227# 0.0172f
C1212 w_n1594_34626# a_1500_33490# 0.0023f
C1213 a_1500_33490# a_1500_34726# 0.0105f
C1214 a_n1500_59349# w_n1594_58110# 0.0172f
C1215 a_1500_16186# a_1500_14950# 0.0105f
C1216 a_n1500_14853# a_n1558_14950# 0.217f
C1217 w_n1594_37098# a_1500_37198# 0.0187f
C1218 a_n1500_n53127# a_n1500_n54363# 3.11f
C1219 a_n1500_n14811# a_n1500_n16047# 3.11f
C1220 a_n1500_30921# w_n1594_32154# 0.0172f
C1221 a_1500_n23366# a_1500_n24602# 0.0105f
C1222 w_n1594_n24702# a_1500_n25838# 0.0023f
C1223 w_n1594_18# a_n1558_1354# 0.0023f
C1224 a_n1500_n24699# a_n1558_n24602# 0.217f
C1225 w_n1594_n6162# a_n1500_n7395# 0.0172f
C1226 a_n1500_42045# a_n1558_42142# 0.217f
C1227 a_1500_52030# w_n1594_53166# 0.0023f
C1228 a_1500_43378# a_1500_42142# 0.0105f
C1229 a_n1558_1354# a_n1558_118# 0.0105f
C1230 w_n1594_35862# a_n1500_35865# 1.65f
C1231 w_n1594_49458# a_n1500_48225# 0.0172f
C1232 a_n1500_35865# a_1500_35962# 0.217f
C1233 a_1500_n41906# w_n1594_n42006# 0.0187f
C1234 w_n1594_51930# a_n1500_51933# 1.65f
C1235 a_1500_n6062# a_1500_n7298# 0.0105f
C1236 a_n1500_n7395# a_n1558_n7298# 0.217f
C1237 a_n1558_n12242# w_n1594_n13578# 0.0023f
C1238 a_n1558_n38198# w_n1594_n37062# 0.0023f
C1239 a_n1558_6298# a_n1558_5062# 0.0105f
C1240 a_n1500_28449# a_n1500_27213# 3.11f
C1241 a_n1500_n17283# w_n1594_n18522# 0.0172f
C1242 a_1500_n8534# w_n1594_n8634# 0.0187f
C1243 a_n1500_n34587# w_n1594_n35826# 0.0172f
C1244 a_n1500_21033# a_n1500_19797# 3.11f
C1245 w_n1594_n60546# a_1500_n60446# 0.0187f
C1246 w_n1594_n7398# a_n1558_n6062# 0.0023f
C1247 a_n1558_n46850# a_n1558_n48086# 0.0105f
C1248 w_n1594_n27174# a_1500_n25838# 0.0023f
C1249 a_1500_47086# w_n1594_45750# 0.0023f
C1250 w_n1594_27210# a_n1558_27310# 0.0187f
C1251 a_1500_n49322# w_n1594_n48186# 0.0023f
C1252 a_n1558_n45614# w_n1594_n46950# 0.0023f
C1253 w_n1594_29682# a_1500_31018# 0.0023f
C1254 a_1500_32254# w_n1594_33390# 0.0023f
C1255 a_n1500_n34587# a_1500_n34490# 0.217f
C1256 w_n1594_42042# a_n1558_43378# 0.0023f
C1257 a_n1500_8673# w_n1594_8670# 1.65f
C1258 w_n1594_n4926# a_1500_n4826# 0.0187f
C1259 a_n1500_n59307# a_n1500_n60543# 3.11f
C1260 a_n1500_n1215# a_n1500_n2451# 3.11f
C1261 a_n1500_n19755# w_n1594_n20994# 0.0172f
C1262 w_n1594_13614# a_n1500_13617# 1.65f
C1263 a_1500_12478# a_1500_11242# 0.0105f
C1264 a_n1500_11145# a_n1558_11242# 0.217f
C1265 a_n1500_11145# w_n1594_11142# 1.65f
C1266 w_n1594_38334# a_n1558_38434# 0.0187f
C1267 a_n1500_51933# a_1500_52030# 0.217f
C1268 w_n1594_n32118# a_n1558_n32018# 0.0187f
C1269 a_1500_n54266# w_n1594_n53130# 0.0023f
C1270 a_n1500_n43239# a_n1500_n44475# 3.11f
C1271 a_n1558_n50558# w_n1594_n51894# 0.0023f
C1272 w_n1594_16086# a_1500_16186# 0.0187f
C1273 a_n1558_n33254# w_n1594_n32118# 0.0023f
C1274 a_n1558_n20894# w_n1594_n19758# 0.0023f
C1275 a_n1500_7437# w_n1594_7434# 1.65f
C1276 a_1500_49558# a_1500_48322# 0.0105f
C1277 a_1500_n35726# w_n1594_n34590# 0.0023f
C1278 w_n1594_39570# a_n1500_38337# 0.0172f
C1279 a_n1500_n50655# a_1500_n50558# 0.217f
C1280 w_n1594_n58074# a_n1500_n59307# 0.0172f
C1281 a_n1500_n20991# a_1500_n20894# 0.217f
C1282 w_n1594_17322# a_n1558_16186# 0.0023f
C1283 a_n1500_n12339# a_1500_n12242# 0.217f
C1284 w_n1594_n25938# a_1500_n24602# 0.0023f
C1285 w_n1594_n22230# a_n1500_n22227# 1.65f
C1286 a_1500_n55502# a_1500_n56738# 0.0105f
C1287 a_n1558_44614# w_n1594_43278# 0.0023f
C1288 w_n1594_44514# a_n1558_43378# 0.0023f
C1289 a_n1558_n36962# a_n1558_n38198# 0.0105f
C1290 w_n1594_n55602# a_n1500_n56835# 0.0172f
C1291 a_n1500_38337# a_n1558_38434# 0.217f
C1292 a_1500_39670# a_1500_38434# 0.0105f
C1293 a_n1558_13714# w_n1594_12378# 0.0023f
C1294 a_n1558_7534# w_n1594_6198# 0.0023f
C1295 a_1500_n40670# w_n1594_n39534# 0.0023f
C1296 a_n1558_n36962# w_n1594_n38298# 0.0023f
C1297 a_n1500_55641# w_n1594_54402# 0.0172f
C1298 a_1500_55738# w_n1594_56874# 0.0023f
C1299 a_n1558_55738# w_n1594_55638# 0.0187f
C1300 a_n1558_3826# w_n1594_4962# 0.0023f
C1301 a_n1500_30921# a_1500_31018# 0.217f
C1302 a_n1500_23505# a_1500_23602# 0.217f
C1303 a_n1500_n30879# a_n1558_n30782# 0.217f
C1304 a_1500_n29546# a_1500_n30782# 0.0105f
C1305 a_n1558_49558# a_n1558_48322# 0.0105f
C1306 w_n1594_n29646# a_1500_n29546# 0.0187f
C1307 a_1500_n48086# w_n1594_n49422# 0.0023f
C1308 w_n1594_n1218# a_1500_n1118# 0.0187f
C1309 a_n1558_40906# a_n1558_39670# 0.0105f
C1310 a_n1500_55641# a_n1558_55738# 0.217f
C1311 a_1500_56974# a_1500_55738# 0.0105f
C1312 w_n1594_46986# a_n1500_46989# 1.65f
C1313 w_n1594_22266# a_1500_23602# 0.0023f
C1314 w_n1594_n23466# a_1500_n22130# 0.0023f
C1315 a_n1500_14853# a_n1500_13617# 3.11f
C1316 a_n1500_32157# a_n1500_33393# 3.11f
C1317 a_n1558_n13478# w_n1594_n14814# 0.0023f
C1318 w_n1594_37098# a_n1558_35962# 0.0023f
C1319 a_n1558_n9770# w_n1594_n11106# 0.0023f
C1320 a_n1558_n53030# a_n1558_n54266# 0.0105f
C1321 a_n1558_n14714# a_n1558_n15950# 0.0105f
C1322 a_n1558_39670# w_n1594_40806# 0.0023f
C1323 a_1500_31018# w_n1594_32154# 0.0023f
C1324 w_n1594_18# a_n1500_21# 1.65f
C1325 a_n1500_n24699# a_n1500_n25935# 3.11f
C1326 w_n1594_n6162# a_1500_n7298# 0.0023f
C1327 a_n1500_4965# w_n1594_3726# 0.0172f
C1328 a_n1558_32254# w_n1594_30918# 0.0023f
C1329 a_n1500_42045# a_n1500_40809# 3.11f
C1330 a_n1500_21# a_n1558_118# 0.217f
C1331 a_1500_1354# a_1500_118# 0.0105f
C1332 a_n1500_n45711# w_n1594_n44478# 0.0172f
C1333 a_n1500_n40767# a_1500_n40670# 0.217f
C1334 w_n1594_35862# a_1500_35962# 0.0187f
C1335 a_n1558_n43142# w_n1594_n42006# 0.0023f
C1336 a_n1500_n7395# a_n1500_n8631# 3.11f
C1337 w_n1594_28446# a_n1558_29782# 0.0023f
C1338 a_n1500_n39531# w_n1594_n40770# 0.0172f
C1339 w_n1594_51930# a_1500_52030# 0.0187f
C1340 a_n1500_n13575# w_n1594_n13578# 1.65f
C1341 a_n1500_4965# a_n1558_5062# 0.217f
C1342 a_n1558_28546# a_n1558_27310# 0.0105f
C1343 w_n1594_46986# a_n1558_48322# 0.0023f
C1344 a_1500_6298# a_1500_5062# 0.0105f
C1345 a_n1558_21130# a_n1558_19894# 0.0105f
C1346 a_1500_n34490# w_n1594_n35826# 0.0023f
C1347 a_1500_n17186# w_n1594_n18522# 0.0023f
C1348 w_n1594_n60546# a_n1558_n61682# 0.0023f
C1349 w_n1594_n59310# a_n1500_n58071# 0.0172f
C1350 w_n1594_n7398# a_n1500_n7395# 1.65f
C1351 a_n1500_n48183# a_n1558_n48086# 0.217f
C1352 w_n1594_n27174# a_n1558_n27074# 0.0187f
C1353 a_1500_n46850# a_1500_n48086# 0.0105f
C1354 a_n1558_n14714# w_n1594_n16050# 0.0023f
C1355 a_n1500_n9867# a_n1558_n9770# 0.217f
C1356 a_n1558_60682# a_n1558_59446# 0.0105f
C1357 a_n1500_n45711# a_1500_n45614# 0.217f
C1358 w_n1594_18558# a_n1558_19894# 0.0023f
C1359 a_n1558_45850# w_n1594_45750# 0.0187f
C1360 w_n1594_27210# a_n1500_25977# 0.0172f
C1361 a_n1500_n46947# w_n1594_n46950# 1.65f
C1362 a_n1500_n44475# w_n1594_n45714# 0.0172f
C1363 w_n1594_29682# a_n1558_29782# 0.0187f
C1364 w_n1594_n56838# a_n1500_n55599# 0.0172f
C1365 w_n1594_42042# a_n1500_42045# 1.65f
C1366 a_1500_8770# w_n1594_8670# 0.0187f
C1367 a_n1558_n59210# a_n1558_n60446# 0.0105f
C1368 w_n1594_n4926# a_n1558_n6062# 0.0023f
C1369 a_n1558_n1118# a_n1558_n2354# 0.0105f
C1370 w_n1594_23502# a_1500_24838# 0.0023f
C1371 w_n1594_n19758# a_1500_n20894# 0.0023f
C1372 a_1500_n19658# w_n1594_n20994# 0.0023f
C1373 a_n1500_n18519# a_1500_n18422# 0.217f
C1374 a_n1500_11145# a_n1500_9909# 3.11f
C1375 a_1500_11242# w_n1594_11142# 0.0187f
C1376 w_n1594_38334# a_n1500_37101# 0.0172f
C1377 w_n1594_n32118# a_n1500_n33351# 0.0172f
C1378 a_n1500_n51891# w_n1594_n51894# 1.65f
C1379 a_n1558_n43142# a_n1558_n44378# 0.0105f
C1380 a_n1558_58210# w_n1594_58110# 0.0187f
C1381 w_n1594_16086# a_n1558_14950# 0.0023f
C1382 w_n1594_n33354# a_n1500_n32115# 0.0172f
C1383 a_n1558_59446# w_n1594_59346# 0.0187f
C1384 a_1500_7534# w_n1594_7434# 0.0187f
C1385 a_n1500_48225# a_n1500_46989# 3.11f
C1386 w_n1594_39570# a_1500_38434# 0.0023f
C1387 a_n1500_17325# a_1500_17422# 0.217f
C1388 w_n1594_n58074# a_1500_n59210# 0.0023f
C1389 w_n1594_21030# a_n1500_22269# 0.0172f
C1390 w_n1594_n25938# a_n1558_n25838# 0.0187f
C1391 a_1500_n61682# VSUBS 0.638f
C1392 a_n1558_n61682# VSUBS 0.638f
C1393 a_n1500_n61779# VSUBS 5.03f
C1394 a_1500_n60446# VSUBS 0.625f
C1395 a_n1558_n60446# VSUBS 0.625f
C1396 a_n1500_n60543# VSUBS 3.31f
C1397 a_1500_n59210# VSUBS 0.625f
C1398 a_n1558_n59210# VSUBS 0.625f
C1399 a_n1500_n59307# VSUBS 3.31f
C1400 a_1500_n57974# VSUBS 0.625f
C1401 a_n1558_n57974# VSUBS 0.625f
C1402 a_n1500_n58071# VSUBS 3.31f
C1403 a_1500_n56738# VSUBS 0.625f
C1404 a_n1558_n56738# VSUBS 0.625f
C1405 a_n1500_n56835# VSUBS 3.31f
C1406 a_1500_n55502# VSUBS 0.625f
C1407 a_n1558_n55502# VSUBS 0.625f
C1408 a_n1500_n55599# VSUBS 3.31f
C1409 a_1500_n54266# VSUBS 0.625f
C1410 a_n1558_n54266# VSUBS 0.625f
C1411 a_n1500_n54363# VSUBS 3.31f
C1412 a_1500_n53030# VSUBS 0.625f
C1413 a_n1558_n53030# VSUBS 0.625f
C1414 a_n1500_n53127# VSUBS 3.31f
C1415 a_1500_n51794# VSUBS 0.625f
C1416 a_n1558_n51794# VSUBS 0.625f
C1417 a_n1500_n51891# VSUBS 3.31f
C1418 a_1500_n50558# VSUBS 0.625f
C1419 a_n1558_n50558# VSUBS 0.625f
C1420 a_n1500_n50655# VSUBS 3.31f
C1421 a_1500_n49322# VSUBS 0.625f
C1422 a_n1558_n49322# VSUBS 0.625f
C1423 a_n1500_n49419# VSUBS 3.31f
C1424 a_1500_n48086# VSUBS 0.625f
C1425 a_n1558_n48086# VSUBS 0.625f
C1426 a_n1500_n48183# VSUBS 3.31f
C1427 a_1500_n46850# VSUBS 0.625f
C1428 a_n1558_n46850# VSUBS 0.625f
C1429 a_n1500_n46947# VSUBS 3.31f
C1430 a_1500_n45614# VSUBS 0.625f
C1431 a_n1558_n45614# VSUBS 0.625f
C1432 a_n1500_n45711# VSUBS 3.31f
C1433 a_1500_n44378# VSUBS 0.625f
C1434 a_n1558_n44378# VSUBS 0.625f
C1435 a_n1500_n44475# VSUBS 3.31f
C1436 a_1500_n43142# VSUBS 0.625f
C1437 a_n1558_n43142# VSUBS 0.625f
C1438 a_n1500_n43239# VSUBS 3.31f
C1439 a_1500_n41906# VSUBS 0.625f
C1440 a_n1558_n41906# VSUBS 0.625f
C1441 a_n1500_n42003# VSUBS 3.31f
C1442 a_1500_n40670# VSUBS 0.625f
C1443 a_n1558_n40670# VSUBS 0.625f
C1444 a_n1500_n40767# VSUBS 3.31f
C1445 a_1500_n39434# VSUBS 0.625f
C1446 a_n1558_n39434# VSUBS 0.625f
C1447 a_n1500_n39531# VSUBS 3.31f
C1448 a_1500_n38198# VSUBS 0.625f
C1449 a_n1558_n38198# VSUBS 0.625f
C1450 a_n1500_n38295# VSUBS 3.31f
C1451 a_1500_n36962# VSUBS 0.625f
C1452 a_n1558_n36962# VSUBS 0.625f
C1453 a_n1500_n37059# VSUBS 3.31f
C1454 a_1500_n35726# VSUBS 0.625f
C1455 a_n1558_n35726# VSUBS 0.625f
C1456 a_n1500_n35823# VSUBS 3.31f
C1457 a_1500_n34490# VSUBS 0.625f
C1458 a_n1558_n34490# VSUBS 0.625f
C1459 a_n1500_n34587# VSUBS 3.31f
C1460 a_1500_n33254# VSUBS 0.625f
C1461 a_n1558_n33254# VSUBS 0.625f
C1462 a_n1500_n33351# VSUBS 3.31f
C1463 a_1500_n32018# VSUBS 0.625f
C1464 a_n1558_n32018# VSUBS 0.625f
C1465 a_n1500_n32115# VSUBS 3.31f
C1466 a_1500_n30782# VSUBS 0.625f
C1467 a_n1558_n30782# VSUBS 0.625f
C1468 a_n1500_n30879# VSUBS 3.31f
C1469 a_1500_n29546# VSUBS 0.625f
C1470 a_n1558_n29546# VSUBS 0.625f
C1471 a_n1500_n29643# VSUBS 3.31f
C1472 a_1500_n28310# VSUBS 0.625f
C1473 a_n1558_n28310# VSUBS 0.625f
C1474 a_n1500_n28407# VSUBS 3.31f
C1475 a_1500_n27074# VSUBS 0.625f
C1476 a_n1558_n27074# VSUBS 0.625f
C1477 a_n1500_n27171# VSUBS 3.31f
C1478 a_1500_n25838# VSUBS 0.625f
C1479 a_n1558_n25838# VSUBS 0.625f
C1480 a_n1500_n25935# VSUBS 3.31f
C1481 a_1500_n24602# VSUBS 0.625f
C1482 a_n1558_n24602# VSUBS 0.625f
C1483 a_n1500_n24699# VSUBS 3.31f
C1484 a_1500_n23366# VSUBS 0.625f
C1485 a_n1558_n23366# VSUBS 0.625f
C1486 a_n1500_n23463# VSUBS 3.31f
C1487 a_1500_n22130# VSUBS 0.625f
C1488 a_n1558_n22130# VSUBS 0.625f
C1489 a_n1500_n22227# VSUBS 3.31f
C1490 a_1500_n20894# VSUBS 0.625f
C1491 a_n1558_n20894# VSUBS 0.625f
C1492 a_n1500_n20991# VSUBS 3.31f
C1493 a_1500_n19658# VSUBS 0.625f
C1494 a_n1558_n19658# VSUBS 0.625f
C1495 a_n1500_n19755# VSUBS 3.31f
C1496 a_1500_n18422# VSUBS 0.625f
C1497 a_n1558_n18422# VSUBS 0.625f
C1498 a_n1500_n18519# VSUBS 3.31f
C1499 a_1500_n17186# VSUBS 0.625f
C1500 a_n1558_n17186# VSUBS 0.625f
C1501 a_n1500_n17283# VSUBS 3.31f
C1502 a_1500_n15950# VSUBS 0.625f
C1503 a_n1558_n15950# VSUBS 0.625f
C1504 a_n1500_n16047# VSUBS 3.31f
C1505 a_1500_n14714# VSUBS 0.625f
C1506 a_n1558_n14714# VSUBS 0.625f
C1507 a_n1500_n14811# VSUBS 3.31f
C1508 a_1500_n13478# VSUBS 0.625f
C1509 a_n1558_n13478# VSUBS 0.625f
C1510 a_n1500_n13575# VSUBS 3.31f
C1511 a_1500_n12242# VSUBS 0.625f
C1512 a_n1558_n12242# VSUBS 0.625f
C1513 a_n1500_n12339# VSUBS 3.31f
C1514 a_1500_n11006# VSUBS 0.625f
C1515 a_n1558_n11006# VSUBS 0.625f
C1516 a_n1500_n11103# VSUBS 3.31f
C1517 a_1500_n9770# VSUBS 0.625f
C1518 a_n1558_n9770# VSUBS 0.625f
C1519 a_n1500_n9867# VSUBS 3.31f
C1520 a_1500_n8534# VSUBS 0.625f
C1521 a_n1558_n8534# VSUBS 0.625f
C1522 a_n1500_n8631# VSUBS 3.31f
C1523 a_1500_n7298# VSUBS 0.625f
C1524 a_n1558_n7298# VSUBS 0.625f
C1525 a_n1500_n7395# VSUBS 3.31f
C1526 a_1500_n6062# VSUBS 0.625f
C1527 a_n1558_n6062# VSUBS 0.625f
C1528 a_n1500_n6159# VSUBS 3.31f
C1529 a_1500_n4826# VSUBS 0.625f
C1530 a_n1558_n4826# VSUBS 0.625f
C1531 a_n1500_n4923# VSUBS 3.31f
C1532 a_1500_n3590# VSUBS 0.625f
C1533 a_n1558_n3590# VSUBS 0.625f
C1534 a_n1500_n3687# VSUBS 3.31f
C1535 a_1500_n2354# VSUBS 0.625f
C1536 a_n1558_n2354# VSUBS 0.625f
C1537 a_n1500_n2451# VSUBS 3.31f
C1538 a_1500_n1118# VSUBS 0.625f
C1539 a_n1558_n1118# VSUBS 0.625f
C1540 a_n1500_n1215# VSUBS 3.31f
C1541 a_1500_118# VSUBS 0.625f
C1542 a_n1558_118# VSUBS 0.625f
C1543 a_n1500_21# VSUBS 3.31f
C1544 a_1500_1354# VSUBS 0.625f
C1545 a_n1558_1354# VSUBS 0.625f
C1546 a_n1500_1257# VSUBS 3.31f
C1547 a_1500_2590# VSUBS 0.625f
C1548 a_n1558_2590# VSUBS 0.625f
C1549 a_n1500_2493# VSUBS 3.31f
C1550 a_1500_3826# VSUBS 0.625f
C1551 a_n1558_3826# VSUBS 0.625f
C1552 a_n1500_3729# VSUBS 3.31f
C1553 a_1500_5062# VSUBS 0.625f
C1554 a_n1558_5062# VSUBS 0.625f
C1555 a_n1500_4965# VSUBS 3.31f
C1556 a_1500_6298# VSUBS 0.625f
C1557 a_n1558_6298# VSUBS 0.625f
C1558 a_n1500_6201# VSUBS 3.31f
C1559 a_1500_7534# VSUBS 0.625f
C1560 a_n1558_7534# VSUBS 0.625f
C1561 a_n1500_7437# VSUBS 3.31f
C1562 a_1500_8770# VSUBS 0.625f
C1563 a_n1558_8770# VSUBS 0.625f
C1564 a_n1500_8673# VSUBS 3.31f
C1565 a_1500_10006# VSUBS 0.625f
C1566 a_n1558_10006# VSUBS 0.625f
C1567 a_n1500_9909# VSUBS 3.31f
C1568 a_1500_11242# VSUBS 0.625f
C1569 a_n1558_11242# VSUBS 0.625f
C1570 a_n1500_11145# VSUBS 3.31f
C1571 a_1500_12478# VSUBS 0.625f
C1572 a_n1558_12478# VSUBS 0.625f
C1573 a_n1500_12381# VSUBS 3.31f
C1574 a_1500_13714# VSUBS 0.625f
C1575 a_n1558_13714# VSUBS 0.625f
C1576 a_n1500_13617# VSUBS 3.31f
C1577 a_1500_14950# VSUBS 0.625f
C1578 a_n1558_14950# VSUBS 0.625f
C1579 a_n1500_14853# VSUBS 3.31f
C1580 a_1500_16186# VSUBS 0.625f
C1581 a_n1558_16186# VSUBS 0.625f
C1582 a_n1500_16089# VSUBS 3.31f
C1583 a_1500_17422# VSUBS 0.625f
C1584 a_n1558_17422# VSUBS 0.625f
C1585 a_n1500_17325# VSUBS 3.31f
C1586 a_1500_18658# VSUBS 0.625f
C1587 a_n1558_18658# VSUBS 0.625f
C1588 a_n1500_18561# VSUBS 3.31f
C1589 a_1500_19894# VSUBS 0.625f
C1590 a_n1558_19894# VSUBS 0.625f
C1591 a_n1500_19797# VSUBS 3.31f
C1592 a_1500_21130# VSUBS 0.625f
C1593 a_n1558_21130# VSUBS 0.625f
C1594 a_n1500_21033# VSUBS 3.31f
C1595 a_1500_22366# VSUBS 0.625f
C1596 a_n1558_22366# VSUBS 0.625f
C1597 a_n1500_22269# VSUBS 3.31f
C1598 a_1500_23602# VSUBS 0.625f
C1599 a_n1558_23602# VSUBS 0.625f
C1600 a_n1500_23505# VSUBS 3.31f
C1601 a_1500_24838# VSUBS 0.625f
C1602 a_n1558_24838# VSUBS 0.625f
C1603 a_n1500_24741# VSUBS 3.31f
C1604 a_1500_26074# VSUBS 0.625f
C1605 a_n1558_26074# VSUBS 0.625f
C1606 a_n1500_25977# VSUBS 3.31f
C1607 a_1500_27310# VSUBS 0.625f
C1608 a_n1558_27310# VSUBS 0.625f
C1609 a_n1500_27213# VSUBS 3.31f
C1610 a_1500_28546# VSUBS 0.625f
C1611 a_n1558_28546# VSUBS 0.625f
C1612 a_n1500_28449# VSUBS 3.31f
C1613 a_1500_29782# VSUBS 0.625f
C1614 a_n1558_29782# VSUBS 0.625f
C1615 a_n1500_29685# VSUBS 3.31f
C1616 a_1500_31018# VSUBS 0.625f
C1617 a_n1558_31018# VSUBS 0.625f
C1618 a_n1500_30921# VSUBS 3.31f
C1619 a_1500_32254# VSUBS 0.625f
C1620 a_n1558_32254# VSUBS 0.625f
C1621 a_n1500_32157# VSUBS 3.31f
C1622 a_1500_33490# VSUBS 0.625f
C1623 a_n1558_33490# VSUBS 0.625f
C1624 a_n1500_33393# VSUBS 3.31f
C1625 a_1500_34726# VSUBS 0.625f
C1626 a_n1558_34726# VSUBS 0.625f
C1627 a_n1500_34629# VSUBS 3.31f
C1628 a_1500_35962# VSUBS 0.625f
C1629 a_n1558_35962# VSUBS 0.625f
C1630 a_n1500_35865# VSUBS 3.31f
C1631 a_1500_37198# VSUBS 0.625f
C1632 a_n1558_37198# VSUBS 0.625f
C1633 a_n1500_37101# VSUBS 3.31f
C1634 a_1500_38434# VSUBS 0.625f
C1635 a_n1558_38434# VSUBS 0.625f
C1636 a_n1500_38337# VSUBS 3.31f
C1637 a_1500_39670# VSUBS 0.625f
C1638 a_n1558_39670# VSUBS 0.625f
C1639 a_n1500_39573# VSUBS 3.31f
C1640 a_1500_40906# VSUBS 0.625f
C1641 a_n1558_40906# VSUBS 0.625f
C1642 a_n1500_40809# VSUBS 3.31f
C1643 a_1500_42142# VSUBS 0.625f
C1644 a_n1558_42142# VSUBS 0.625f
C1645 a_n1500_42045# VSUBS 3.31f
C1646 a_1500_43378# VSUBS 0.625f
C1647 a_n1558_43378# VSUBS 0.625f
C1648 a_n1500_43281# VSUBS 3.31f
C1649 a_1500_44614# VSUBS 0.625f
C1650 a_n1558_44614# VSUBS 0.625f
C1651 a_n1500_44517# VSUBS 3.31f
C1652 a_1500_45850# VSUBS 0.625f
C1653 a_n1558_45850# VSUBS 0.625f
C1654 a_n1500_45753# VSUBS 3.31f
C1655 a_1500_47086# VSUBS 0.625f
C1656 a_n1558_47086# VSUBS 0.625f
C1657 a_n1500_46989# VSUBS 3.31f
C1658 a_1500_48322# VSUBS 0.625f
C1659 a_n1558_48322# VSUBS 0.625f
C1660 a_n1500_48225# VSUBS 3.31f
C1661 a_1500_49558# VSUBS 0.625f
C1662 a_n1558_49558# VSUBS 0.625f
C1663 a_n1500_49461# VSUBS 3.31f
C1664 a_1500_50794# VSUBS 0.625f
C1665 a_n1558_50794# VSUBS 0.625f
C1666 a_n1500_50697# VSUBS 3.31f
C1667 a_1500_52030# VSUBS 0.625f
C1668 a_n1558_52030# VSUBS 0.625f
C1669 a_n1500_51933# VSUBS 3.31f
C1670 a_1500_53266# VSUBS 0.625f
C1671 a_n1558_53266# VSUBS 0.625f
C1672 a_n1500_53169# VSUBS 3.31f
C1673 a_1500_54502# VSUBS 0.625f
C1674 a_n1558_54502# VSUBS 0.625f
C1675 a_n1500_54405# VSUBS 3.31f
C1676 a_1500_55738# VSUBS 0.625f
C1677 a_n1558_55738# VSUBS 0.625f
C1678 a_n1500_55641# VSUBS 3.31f
C1679 a_1500_56974# VSUBS 0.625f
C1680 a_n1558_56974# VSUBS 0.625f
C1681 a_n1500_56877# VSUBS 3.31f
C1682 a_1500_58210# VSUBS 0.625f
C1683 a_n1558_58210# VSUBS 0.625f
C1684 a_n1500_58113# VSUBS 3.31f
C1685 a_1500_59446# VSUBS 0.625f
C1686 a_n1558_59446# VSUBS 0.625f
C1687 a_n1500_59349# VSUBS 3.31f
C1688 a_1500_60682# VSUBS 0.638f
C1689 a_n1558_60682# VSUBS 0.638f
C1690 a_n1500_60585# VSUBS 5.03f
C1691 w_n1594_n61782# VSUBS 11.5f
C1692 w_n1594_n60546# VSUBS 11.5f
C1693 w_n1594_n59310# VSUBS 11.5f
C1694 w_n1594_n58074# VSUBS 11.5f
C1695 w_n1594_n56838# VSUBS 11.5f
C1696 w_n1594_n55602# VSUBS 11.5f
C1697 w_n1594_n54366# VSUBS 11.5f
C1698 w_n1594_n53130# VSUBS 11.5f
C1699 w_n1594_n51894# VSUBS 11.5f
C1700 w_n1594_n50658# VSUBS 11.5f
C1701 w_n1594_n49422# VSUBS 11.5f
C1702 w_n1594_n48186# VSUBS 11.5f
C1703 w_n1594_n46950# VSUBS 11.5f
C1704 w_n1594_n45714# VSUBS 11.5f
C1705 w_n1594_n44478# VSUBS 11.5f
C1706 w_n1594_n43242# VSUBS 11.5f
C1707 w_n1594_n42006# VSUBS 11.5f
C1708 w_n1594_n40770# VSUBS 11.5f
C1709 w_n1594_n39534# VSUBS 11.5f
C1710 w_n1594_n38298# VSUBS 11.5f
C1711 w_n1594_n37062# VSUBS 11.5f
C1712 w_n1594_n35826# VSUBS 11.5f
C1713 w_n1594_n34590# VSUBS 11.5f
C1714 w_n1594_n33354# VSUBS 11.5f
C1715 w_n1594_n32118# VSUBS 11.5f
C1716 w_n1594_n30882# VSUBS 11.5f
C1717 w_n1594_n29646# VSUBS 11.5f
C1718 w_n1594_n28410# VSUBS 11.5f
C1719 w_n1594_n27174# VSUBS 11.5f
C1720 w_n1594_n25938# VSUBS 11.5f
C1721 w_n1594_n24702# VSUBS 11.5f
C1722 w_n1594_n23466# VSUBS 11.5f
C1723 w_n1594_n22230# VSUBS 11.5f
C1724 w_n1594_n20994# VSUBS 11.5f
C1725 w_n1594_n19758# VSUBS 11.5f
C1726 w_n1594_n18522# VSUBS 11.5f
C1727 w_n1594_n17286# VSUBS 11.5f
C1728 w_n1594_n16050# VSUBS 11.5f
C1729 w_n1594_n14814# VSUBS 11.5f
C1730 w_n1594_n13578# VSUBS 11.5f
C1731 w_n1594_n12342# VSUBS 11.5f
C1732 w_n1594_n11106# VSUBS 11.5f
C1733 w_n1594_n9870# VSUBS 11.5f
C1734 w_n1594_n8634# VSUBS 11.5f
C1735 w_n1594_n7398# VSUBS 11.5f
C1736 w_n1594_n6162# VSUBS 11.5f
C1737 w_n1594_n4926# VSUBS 11.5f
C1738 w_n1594_n3690# VSUBS 11.5f
C1739 w_n1594_n2454# VSUBS 11.5f
C1740 w_n1594_n1218# VSUBS 11.5f
C1741 w_n1594_18# VSUBS 11.5f
C1742 w_n1594_1254# VSUBS 11.5f
C1743 w_n1594_2490# VSUBS 11.5f
C1744 w_n1594_3726# VSUBS 11.5f
C1745 w_n1594_4962# VSUBS 11.5f
C1746 w_n1594_6198# VSUBS 11.5f
C1747 w_n1594_7434# VSUBS 11.5f
C1748 w_n1594_8670# VSUBS 11.5f
C1749 w_n1594_9906# VSUBS 11.5f
C1750 w_n1594_11142# VSUBS 11.5f
C1751 w_n1594_12378# VSUBS 11.5f
C1752 w_n1594_13614# VSUBS 11.5f
C1753 w_n1594_14850# VSUBS 11.5f
C1754 w_n1594_16086# VSUBS 11.5f
C1755 w_n1594_17322# VSUBS 11.5f
C1756 w_n1594_18558# VSUBS 11.5f
C1757 w_n1594_19794# VSUBS 11.5f
C1758 w_n1594_21030# VSUBS 11.5f
C1759 w_n1594_22266# VSUBS 11.5f
C1760 w_n1594_23502# VSUBS 11.5f
C1761 w_n1594_24738# VSUBS 11.5f
C1762 w_n1594_25974# VSUBS 11.5f
C1763 w_n1594_27210# VSUBS 11.5f
C1764 w_n1594_28446# VSUBS 11.5f
C1765 w_n1594_29682# VSUBS 11.5f
C1766 w_n1594_30918# VSUBS 11.5f
C1767 w_n1594_32154# VSUBS 11.5f
C1768 w_n1594_33390# VSUBS 11.5f
C1769 w_n1594_34626# VSUBS 11.5f
C1770 w_n1594_35862# VSUBS 11.5f
C1771 w_n1594_37098# VSUBS 11.5f
C1772 w_n1594_38334# VSUBS 11.5f
C1773 w_n1594_39570# VSUBS 11.5f
C1774 w_n1594_40806# VSUBS 11.5f
C1775 w_n1594_42042# VSUBS 11.5f
C1776 w_n1594_43278# VSUBS 11.5f
C1777 w_n1594_44514# VSUBS 11.5f
C1778 w_n1594_45750# VSUBS 11.5f
C1779 w_n1594_46986# VSUBS 11.5f
C1780 w_n1594_48222# VSUBS 11.5f
C1781 w_n1594_49458# VSUBS 11.5f
C1782 w_n1594_50694# VSUBS 11.5f
C1783 w_n1594_51930# VSUBS 11.5f
C1784 w_n1594_53166# VSUBS 11.5f
C1785 w_n1594_54402# VSUBS 11.5f
C1786 w_n1594_55638# VSUBS 11.5f
C1787 w_n1594_56874# VSUBS 11.5f
C1788 w_n1594_58110# VSUBS 11.5f
C1789 w_n1594_59346# VSUBS 11.5f
C1790 w_n1594_60582# VSUBS 11.5f
.ends

.subckt sky130_fd_pr__nfet_01v8_WK8VRD a_n500_9156# a_n558_n10244# a_500_n2936# a_500_n5372#
+ a_n500_n1806# a_500_718# a_n500_3066# a_n500_n4242# a_n500_630# a_n500_n6678# a_n558_1936#
+ a_n558_4372# a_n558_n9026# a_n558_n6590# a_500_n500# a_500_6808# a_n500_6720# a_500_9244#
+ a_500_3154# a_500_n7808# a_n500_n9114# a_500_n4154# a_500_n1718# a_n558_n500# a_n500_n3024#
+ a_n558_6808# a_n558_9244# a_n558_n2936# a_n558_3154# a_n500_n10332# a_n558_n5372#
+ a_n558_718# a_n500_n588# a_n500_5502# a_500_8026# a_500_5590# a_n500_7938# a_500_n9026#
+ a_n500_1848# a_500_n6590# a_n500_4284# a_n500_n5460# a_n558_n7808# a_n500_n7896#
+ a_n558_8026# a_n558_n1718# a_n558_5590# a_n558_n4154# a_500_n10244# a_500_1936#
+ a_500_4372# VSUBS
X0 a_500_n10244# a_n500_n10332# a_n558_n10244# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X1 a_500_4372# a_n500_4284# a_n558_4372# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X2 a_500_n6590# a_n500_n6678# a_n558_n6590# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X3 a_500_5590# a_n500_5502# a_n558_5590# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X4 a_500_n1718# a_n500_n1806# a_n558_n1718# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X5 a_500_n2936# a_n500_n3024# a_n558_n2936# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X6 a_500_n4154# a_n500_n4242# a_n558_n4154# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X7 a_500_718# a_n500_630# a_n558_718# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X8 a_500_n5372# a_n500_n5460# a_n558_n5372# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X9 a_500_6808# a_n500_6720# a_n558_6808# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X10 a_500_8026# a_n500_7938# a_n558_8026# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X11 a_500_n500# a_n500_n588# a_n558_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X12 a_500_9244# a_n500_9156# a_n558_9244# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X13 a_500_1936# a_n500_1848# a_n558_1936# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X14 a_500_n7808# a_n500_n7896# a_n558_n7808# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X15 a_500_3154# a_n500_3066# a_n558_3154# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X16 a_500_n9026# a_n500_n9114# a_n558_n9026# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
C0 a_500_6808# a_500_5590# 0.0113f
C1 a_n558_6808# a_n500_6720# 0.204f
C2 a_n500_5502# a_n558_5590# 0.204f
C3 a_n500_n4242# a_n558_n4154# 0.204f
C4 a_n500_n6678# a_n500_n7896# 1.03f
C5 a_n558_n7808# a_n558_n6590# 0.0113f
C6 a_n500_n588# a_n500_630# 1.03f
C7 a_n500_9156# a_n558_9244# 0.204f
C8 a_n500_6720# a_n500_7938# 1.03f
C9 a_500_n500# a_500_n1718# 0.0113f
C10 a_n558_n5372# a_n558_n6590# 0.0113f
C11 a_n500_9156# a_n500_7938# 1.03f
C12 a_n558_9244# a_500_9244# 0.0663f
C13 a_n500_n9114# a_500_n9026# 0.204f
C14 a_n500_n588# a_n558_n500# 0.204f
C15 a_n500_n9114# a_n500_n10332# 1.03f
C16 a_500_6808# a_n500_6720# 0.204f
C17 a_n558_n4154# a_500_n4154# 0.0663f
C18 a_n500_n4242# a_n500_n5460# 1.03f
C19 a_500_718# a_500_n500# 0.0113f
C20 a_n558_5590# a_n558_4372# 0.0113f
C21 a_n558_9244# a_n558_8026# 0.0113f
C22 a_n558_6808# a_n558_8026# 0.0113f
C23 a_n558_n4154# a_n558_n5372# 0.0113f
C24 a_n558_n500# a_500_n500# 0.0663f
C25 a_500_n5372# a_500_n6590# 0.0113f
C26 a_n558_n10244# a_n558_n9026# 0.0113f
C27 a_n500_7938# a_n558_8026# 0.204f
C28 a_500_9244# a_500_8026# 0.0113f
C29 a_n500_n6678# a_n558_n6590# 0.204f
C30 a_n500_3066# a_n558_3154# 0.204f
C31 a_n558_6808# a_n558_5590# 0.0113f
C32 a_500_4372# a_500_5590# 0.0113f
C33 a_n558_8026# a_500_8026# 0.0663f
C34 a_n500_1848# a_500_1936# 0.204f
C35 a_500_n2936# a_n500_n3024# 0.204f
C36 a_n500_n5460# a_n558_n5372# 0.204f
C37 a_n558_n1718# a_500_n1718# 0.0663f
C38 a_n500_n9114# a_n500_n7896# 1.03f
C39 a_500_n2936# a_500_n1718# 0.0113f
C40 a_500_4372# a_n500_4284# 0.204f
C41 a_n558_n2936# a_n558_n4154# 0.0113f
C42 a_500_n5372# a_500_n4154# 0.0113f
C43 a_n500_n588# a_n500_n1806# 1.03f
C44 a_500_n9026# a_500_n10244# 0.0113f
C45 a_n500_n10332# a_500_n10244# 0.204f
C46 a_n500_n4242# a_n500_n3024# 1.03f
C47 a_n558_3154# a_500_3154# 0.0663f
C48 a_500_n5372# a_n558_n5372# 0.0663f
C49 a_n558_n500# a_n558_n1718# 0.0113f
C50 a_n500_n9114# a_n558_n9026# 0.204f
C51 a_500_718# a_n500_630# 0.204f
C52 a_n500_n5460# a_n500_n6678# 1.03f
C53 a_n500_3066# a_n500_4284# 1.03f
C54 a_n558_718# a_n558_1936# 0.0113f
C55 a_n500_3066# a_n500_1848# 1.03f
C56 a_n500_5502# a_500_5590# 0.204f
C57 a_500_n2936# a_500_n4154# 0.0113f
C58 a_n558_5590# a_500_5590# 0.0663f
C59 a_n558_3154# a_n558_4372# 0.0113f
C60 a_n500_9156# a_500_9244# 0.204f
C61 a_500_n7808# a_500_n9026# 0.0113f
C62 a_n558_718# a_n500_630# 0.204f
C63 a_n558_3154# a_n558_1936# 0.0113f
C64 a_n500_5502# a_n500_4284# 1.03f
C65 a_n500_n4242# a_500_n4154# 0.204f
C66 a_500_718# a_n558_718# 0.0663f
C67 a_500_n7808# a_500_n6590# 0.0113f
C68 a_n500_5502# a_n500_6720# 1.03f
C69 a_n558_n500# a_n558_718# 0.0113f
C70 a_n500_n588# a_500_n500# 0.204f
C71 a_500_n9026# a_n558_n9026# 0.0663f
C72 a_500_3154# a_500_1936# 0.0113f
C73 a_n500_n1806# a_n558_n1718# 0.204f
C74 a_n558_n7808# a_n500_n7896# 0.204f
C75 a_n558_n7808# a_500_n7808# 0.0663f
C76 a_n500_4284# a_n558_4372# 0.204f
C77 a_n558_6808# a_500_6808# 0.0663f
C78 a_n558_n2936# a_n558_n1718# 0.0113f
C79 a_n558_n2936# a_500_n2936# 0.0663f
C80 a_n500_7938# a_500_8026# 0.204f
C81 a_n500_n6678# a_500_n6590# 0.204f
C82 a_n500_n3024# a_n500_n1806# 1.03f
C83 a_n500_1848# a_n558_1936# 0.204f
C84 a_500_3154# a_500_4372# 0.0113f
C85 a_n558_n2936# a_n500_n3024# 0.204f
C86 a_n500_n1806# a_500_n1718# 0.204f
C87 a_500_n7808# a_n500_n7896# 0.204f
C88 a_n558_n6590# a_500_n6590# 0.0663f
C89 a_n558_n7808# a_n558_n9026# 0.0113f
C90 a_n558_1936# a_500_1936# 0.0663f
C91 a_n500_1848# a_n500_630# 1.03f
C92 a_n500_n10332# a_n558_n10244# 0.204f
C93 a_500_6808# a_500_8026# 0.0113f
C94 a_n500_3066# a_500_3154# 0.204f
C95 a_500_4372# a_n558_4372# 0.0663f
C96 a_500_n5372# a_n500_n5460# 0.204f
C97 a_n558_n10244# a_500_n10244# 0.0663f
C98 a_500_718# a_500_1936# 0.0113f
C99 a_500_n10244# VSUBS 0.581f
C100 a_n558_n10244# VSUBS 0.581f
C101 a_n500_n10332# VSUBS 2.28f
C102 a_500_n9026# VSUBS 0.571f
C103 a_n558_n9026# VSUBS 0.571f
C104 a_n500_n9114# VSUBS 1.71f
C105 a_500_n7808# VSUBS 0.571f
C106 a_n558_n7808# VSUBS 0.571f
C107 a_n500_n7896# VSUBS 1.71f
C108 a_500_n6590# VSUBS 0.571f
C109 a_n558_n6590# VSUBS 0.571f
C110 a_n500_n6678# VSUBS 1.71f
C111 a_500_n5372# VSUBS 0.571f
C112 a_n558_n5372# VSUBS 0.571f
C113 a_n500_n5460# VSUBS 1.71f
C114 a_500_n4154# VSUBS 0.571f
C115 a_n558_n4154# VSUBS 0.571f
C116 a_n500_n4242# VSUBS 1.71f
C117 a_500_n2936# VSUBS 0.571f
C118 a_n558_n2936# VSUBS 0.571f
C119 a_n500_n3024# VSUBS 1.71f
C120 a_500_n1718# VSUBS 0.571f
C121 a_n558_n1718# VSUBS 0.571f
C122 a_n500_n1806# VSUBS 1.71f
C123 a_500_n500# VSUBS 0.571f
C124 a_n558_n500# VSUBS 0.571f
C125 a_n500_n588# VSUBS 1.71f
C126 a_500_718# VSUBS 0.571f
C127 a_n558_718# VSUBS 0.571f
C128 a_n500_630# VSUBS 1.71f
C129 a_500_1936# VSUBS 0.571f
C130 a_n558_1936# VSUBS 0.571f
C131 a_n500_1848# VSUBS 1.71f
C132 a_500_3154# VSUBS 0.571f
C133 a_n558_3154# VSUBS 0.571f
C134 a_n500_3066# VSUBS 1.71f
C135 a_500_4372# VSUBS 0.571f
C136 a_n558_4372# VSUBS 0.571f
C137 a_n500_4284# VSUBS 1.71f
C138 a_500_5590# VSUBS 0.571f
C139 a_n558_5590# VSUBS 0.571f
C140 a_n500_5502# VSUBS 1.71f
C141 a_500_6808# VSUBS 0.571f
C142 a_n558_6808# VSUBS 0.571f
C143 a_n500_6720# VSUBS 1.71f
C144 a_500_8026# VSUBS 0.571f
C145 a_n558_8026# VSUBS 0.571f
C146 a_n500_7938# VSUBS 1.71f
C147 a_500_9244# VSUBS 0.581f
C148 a_n558_9244# VSUBS 0.581f
C149 a_n500_9156# VSUBS 2.28f
.ends

.subckt sky130_fd_pr__nfet_01v8_AH5E2K a_500_n500# a_n558_n500# a_n500_n588# VSUBS
X0 a_500_n500# a_n500_n588# a_n558_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
C0 a_n500_n588# a_500_n500# 0.204f
C1 a_n500_n588# a_n558_n500# 0.204f
C2 a_n558_n500# a_500_n500# 0.0663f
C3 a_500_n500# VSUBS 0.592f
C4 a_n558_n500# VSUBS 0.592f
C5 a_n500_n588# VSUBS 2.84f
.ends

.subckt sky130_fd_pr__pfet_01v8_C2U9V5 a_n300_n597# a_300_n500# w_n394_n600# a_n358_n500#
+ VSUBS
X0 a_300_n500# a_n300_n597# a_n358_n500# w_n394_n600# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=3
**devattr s=58000,2116 d=58000,2116
C0 w_n394_n600# a_300_n500# 0.0187f
C1 a_n358_n500# a_300_n500# 0.107f
C2 w_n394_n600# a_n358_n500# 0.0187f
C3 a_n300_n597# a_300_n500# 0.184f
C4 w_n394_n600# a_n300_n597# 0.382f
C5 a_n300_n597# a_n358_n500# 0.184f
C6 a_300_n500# VSUBS 0.548f
C7 a_n358_n500# VSUBS 0.548f
C8 a_n300_n597# VSUBS 1.42f
C9 w_n394_n600# VSUBS 2.84f
.ends

.subckt sky130_fd_pr__nfet_01v8_QP5WRD a_500_n2936# a_500_n5372# a_n500_n1806# a_500_718#
+ a_n500_3066# a_n500_n4242# a_n500_630# a_n500_n6678# a_n558_1936# a_n558_4372# a_n558_n9026#
+ a_n558_n6590# a_500_n500# a_500_6808# a_n500_6720# a_500_3154# a_500_n7808# a_n500_n9114#
+ a_500_n4154# a_500_n1718# a_n558_n500# a_n500_n3024# a_n558_6808# a_n558_n2936#
+ a_n558_3154# a_n558_n5372# a_n558_718# a_n500_n588# a_n500_5502# a_500_8026# a_500_5590#
+ a_n500_7938# a_500_n9026# a_n500_1848# a_500_n6590# a_n500_4284# a_n500_n5460# a_n558_n7808#
+ a_n500_n7896# a_n558_8026# a_n558_n1718# a_n558_5590# a_n558_n4154# a_500_1936#
+ a_500_4372# VSUBS
X0 a_500_4372# a_n500_4284# a_n558_4372# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X1 a_500_n6590# a_n500_n6678# a_n558_n6590# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X2 a_500_5590# a_n500_5502# a_n558_5590# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X3 a_500_n1718# a_n500_n1806# a_n558_n1718# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X4 a_500_n2936# a_n500_n3024# a_n558_n2936# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X5 a_500_n4154# a_n500_n4242# a_n558_n4154# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X6 a_500_718# a_n500_630# a_n558_718# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X7 a_500_n5372# a_n500_n5460# a_n558_n5372# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X8 a_500_6808# a_n500_6720# a_n558_6808# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X9 a_500_8026# a_n500_7938# a_n558_8026# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X10 a_500_n500# a_n500_n588# a_n558_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X11 a_500_1936# a_n500_1848# a_n558_1936# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X12 a_500_n7808# a_n500_n7896# a_n558_n7808# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X13 a_500_3154# a_n500_3066# a_n558_3154# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X14 a_500_n9026# a_n500_n9114# a_n558_n9026# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
C0 a_n558_n1718# a_n558_n500# 0.0113f
C1 a_n500_n5460# a_n500_n6678# 1.03f
C2 a_500_n6590# a_n558_n6590# 0.0663f
C3 a_n500_n5460# a_500_n5372# 0.204f
C4 a_500_1936# a_n500_1848# 0.204f
C5 a_n500_n9114# a_n558_n9026# 0.204f
C6 a_500_n7808# a_500_n9026# 0.0113f
C7 a_n500_n3024# a_500_n2936# 0.204f
C8 a_n558_n4154# a_n558_n2936# 0.0113f
C9 a_500_718# a_500_n500# 0.0113f
C10 a_500_3154# a_500_4372# 0.0113f
C11 a_n558_5590# a_n558_4372# 0.0113f
C12 a_n500_7938# a_n500_6720# 1.03f
C13 a_n558_n5372# a_500_n5372# 0.0663f
C14 a_n500_630# a_n500_1848# 1.03f
C15 a_n500_630# a_n558_718# 0.204f
C16 a_n500_n4242# a_n500_n3024# 1.03f
C17 a_500_n500# a_500_n1718# 0.0113f
C18 a_n500_n1806# a_n558_n1718# 0.204f
C19 a_n500_n9114# a_500_n9026# 0.204f
C20 a_n558_n2936# a_500_n2936# 0.0663f
C21 a_n558_8026# a_n558_6808# 0.0113f
C22 a_n500_1848# a_n558_1936# 0.204f
C23 a_n558_718# a_n558_1936# 0.0113f
C24 a_n558_718# a_500_718# 0.0663f
C25 a_n500_n1806# a_500_n1718# 0.204f
C26 a_n558_n7808# a_500_n7808# 0.0663f
C27 a_500_3154# a_n558_3154# 0.0663f
C28 a_n500_4284# a_500_4372# 0.204f
C29 a_500_8026# a_500_6808# 0.0113f
C30 a_n558_n4154# a_n500_n4242# 0.204f
C31 a_500_n6590# a_n500_n6678# 0.204f
C32 a_500_5590# a_500_6808# 0.0113f
C33 a_n500_3066# a_n500_1848# 1.03f
C34 a_500_n6590# a_500_n5372# 0.0113f
C35 a_n558_4372# a_500_4372# 0.0663f
C36 a_n500_n7896# a_n500_n6678# 1.03f
C37 a_n500_n588# a_n558_n500# 0.204f
C38 a_n558_n1718# a_n558_n2936# 0.0113f
C39 a_n500_n6678# a_n558_n6590# 0.204f
C40 a_n558_n4154# a_n558_n5372# 0.0113f
C41 a_n500_n588# a_500_n500# 0.204f
C42 a_n500_6720# a_n558_6808# 0.204f
C43 a_500_1936# a_500_3154# 0.0113f
C44 a_500_n500# a_n558_n500# 0.0663f
C45 a_n500_n5460# a_n500_n4242# 1.03f
C46 a_n558_3154# a_n558_1936# 0.0113f
C47 a_n500_7938# a_500_8026# 0.204f
C48 a_n500_n588# a_n500_n1806# 1.03f
C49 a_n500_4284# a_n500_5502# 1.03f
C50 a_n558_4372# a_n558_3154# 0.0113f
C51 a_n558_6808# a_500_6808# 0.0663f
C52 a_n558_5590# a_500_5590# 0.0663f
C53 a_n500_n5460# a_n558_n5372# 0.204f
C54 a_500_n4154# a_500_n5372# 0.0113f
C55 a_n558_718# a_n558_n500# 0.0113f
C56 a_n500_3066# a_n558_3154# 0.204f
C57 a_500_n1718# a_500_n2936# 0.0113f
C58 a_n500_5502# a_n500_6720# 1.03f
C59 a_n500_n7896# a_n558_n7808# 0.204f
C60 a_500_1936# a_n558_1936# 0.0663f
C61 a_500_1936# a_500_718# 0.0113f
C62 a_n558_n7808# a_n558_n6590# 0.0113f
C63 a_500_3154# a_n500_3066# 0.204f
C64 a_n500_630# a_500_718# 0.204f
C65 a_n558_n9026# a_500_n9026# 0.0663f
C66 a_500_n7808# a_500_n6590# 0.0113f
C67 a_n558_5590# a_n558_6808# 0.0113f
C68 a_n500_4284# a_n558_4372# 0.204f
C69 a_n500_n7896# a_500_n7808# 0.204f
C70 a_500_5590# a_500_4372# 0.0113f
C71 a_n558_n1718# a_500_n1718# 0.0663f
C72 a_n500_n1806# a_n500_n3024# 1.03f
C73 a_n558_n4154# a_500_n4154# 0.0663f
C74 a_n500_4284# a_n500_3066# 1.03f
C75 a_n500_n7896# a_n500_n9114# 1.03f
C76 a_500_n4154# a_500_n2936# 0.0113f
C77 a_n558_n7808# a_n558_n9026# 0.0113f
C78 a_n558_5590# a_n500_5502# 0.204f
C79 a_n558_n5372# a_n558_n6590# 0.0113f
C80 a_500_n4154# a_n500_n4242# 0.204f
C81 a_n500_7938# a_n558_8026# 0.204f
C82 a_500_5590# a_n500_5502# 0.204f
C83 a_n500_6720# a_500_6808# 0.204f
C84 a_n500_630# a_n500_n588# 1.03f
C85 a_n500_n3024# a_n558_n2936# 0.204f
C86 a_n558_8026# a_500_8026# 0.0663f
C87 a_500_n9026# VSUBS 0.581f
C88 a_n558_n9026# VSUBS 0.581f
C89 a_n500_n9114# VSUBS 2.28f
C90 a_500_n7808# VSUBS 0.571f
C91 a_n558_n7808# VSUBS 0.571f
C92 a_n500_n7896# VSUBS 1.71f
C93 a_500_n6590# VSUBS 0.571f
C94 a_n558_n6590# VSUBS 0.571f
C95 a_n500_n6678# VSUBS 1.71f
C96 a_500_n5372# VSUBS 0.571f
C97 a_n558_n5372# VSUBS 0.571f
C98 a_n500_n5460# VSUBS 1.71f
C99 a_500_n4154# VSUBS 0.571f
C100 a_n558_n4154# VSUBS 0.571f
C101 a_n500_n4242# VSUBS 1.71f
C102 a_500_n2936# VSUBS 0.571f
C103 a_n558_n2936# VSUBS 0.571f
C104 a_n500_n3024# VSUBS 1.71f
C105 a_500_n1718# VSUBS 0.571f
C106 a_n558_n1718# VSUBS 0.571f
C107 a_n500_n1806# VSUBS 1.71f
C108 a_500_n500# VSUBS 0.571f
C109 a_n558_n500# VSUBS 0.571f
C110 a_n500_n588# VSUBS 1.71f
C111 a_500_718# VSUBS 0.571f
C112 a_n558_718# VSUBS 0.571f
C113 a_n500_630# VSUBS 1.71f
C114 a_500_1936# VSUBS 0.571f
C115 a_n558_1936# VSUBS 0.571f
C116 a_n500_1848# VSUBS 1.71f
C117 a_500_3154# VSUBS 0.571f
C118 a_n558_3154# VSUBS 0.571f
C119 a_n500_3066# VSUBS 1.71f
C120 a_500_4372# VSUBS 0.571f
C121 a_n558_4372# VSUBS 0.571f
C122 a_n500_4284# VSUBS 1.71f
C123 a_500_5590# VSUBS 0.571f
C124 a_n558_5590# VSUBS 0.571f
C125 a_n500_5502# VSUBS 1.71f
C126 a_500_6808# VSUBS 0.571f
C127 a_n558_6808# VSUBS 0.571f
C128 a_n500_6720# VSUBS 1.71f
C129 a_500_8026# VSUBS 0.581f
C130 a_n558_8026# VSUBS 0.581f
C131 a_n500_7938# VSUBS 2.28f
.ends

.subckt sky130_fd_pr__pfet_01v8_UDM5A5 a_n558_n7916# a_n500_5583# a_500_1972# a_n558_8152#
+ a_n500_8055# a_500_4444# w_n594_3108# w_n594_6816# a_500_n2972# a_500_736# a_500_n5444#
+ a_n500_n597# w_n594_636# a_500_n500# w_n594_n3072# a_n558_1972# w_n594_n6780# w_n594_n600#
+ a_n500_1875# a_n558_4444# w_n594_n9252# a_n500_4347# a_n558_n6680# a_n558_n9152#
+ a_n500_n5541# a_n500_639# a_500_3208# a_n500_n8013# a_500_6916# a_500_n1736# a_n558_n500#
+ a_500_n4208# w_n594_5580# a_500_n7916# w_n594_8052# w_n594_n5544# a_n558_736# a_n558_3208#
+ w_n594_n8016# a_n558_n2972# a_n558_6916# a_n558_n5444# a_n500_n1833# a_n500_6819#
+ a_n500_n4305# w_n594_1872# a_500_5680# a_n500_n3069# w_n594_4344# a_n500_n6777#
+ a_500_8152# w_n594_n1836# a_n500_n9249# a_500_n6680# w_n594_n4308# a_n500_3111#
+ a_500_n9152# a_n558_n1736# a_n558_n4208# a_n558_5680# VSUBS
X0 a_500_1972# a_n500_1875# a_n558_1972# w_n594_1872# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X1 a_500_6916# a_n500_6819# a_n558_6916# w_n594_6816# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X2 a_500_4444# a_n500_4347# a_n558_4444# w_n594_4344# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X3 a_500_n9152# a_n500_n9249# a_n558_n9152# w_n594_n9252# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X4 a_500_3208# a_n500_3111# a_n558_3208# w_n594_3108# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X5 a_500_n2972# a_n500_n3069# a_n558_n2972# w_n594_n3072# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X6 a_500_n7916# a_n500_n8013# a_n558_n7916# w_n594_n8016# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X7 a_500_n5444# a_n500_n5541# a_n558_n5444# w_n594_n5544# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X8 a_500_n500# a_n500_n597# a_n558_n500# w_n594_n600# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X9 a_500_n1736# a_n500_n1833# a_n558_n1736# w_n594_n1836# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X10 a_500_n4208# a_n500_n4305# a_n558_n4208# w_n594_n4308# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X11 a_500_736# a_n500_639# a_n558_736# w_n594_636# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X12 a_500_n6680# a_n500_n6777# a_n558_n6680# w_n594_n6780# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X13 a_500_5680# a_n500_5583# a_n558_5680# w_n594_5580# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X14 a_500_8152# a_n500_8055# a_n558_8152# w_n594_8052# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
C0 a_500_n7916# a_n558_n7916# 0.0663f
C1 w_n594_n6780# a_n558_n7916# 0.0023f
C2 w_n594_3108# a_n500_3111# 0.593f
C3 w_n594_4344# a_n558_3208# 0.0023f
C4 a_n558_n9152# a_n558_n7916# 0.0105f
C5 a_500_5680# a_500_6916# 0.0105f
C6 a_500_n500# a_500_736# 0.0105f
C7 a_n558_3208# a_500_3208# 0.0663f
C8 a_500_n9152# w_n594_n8016# 0.0023f
C9 w_n594_8052# a_n558_6916# 0.0023f
C10 w_n594_6816# a_n558_8152# 0.0023f
C11 a_500_5680# a_500_4444# 0.0105f
C12 a_n500_4347# a_n558_4444# 0.204f
C13 a_500_736# w_n594_636# 0.0187f
C14 a_500_n7916# w_n594_n6780# 0.0023f
C15 w_n594_3108# a_n558_3208# 0.0187f
C16 a_n558_n2972# a_n558_n1736# 0.0105f
C17 a_n500_n1833# a_n558_n1736# 0.204f
C18 a_500_5680# a_n500_5583# 0.204f
C19 w_n594_n5544# a_n500_n5541# 0.593f
C20 a_n558_736# w_n594_636# 0.0187f
C21 a_n558_5680# a_n500_5583# 0.204f
C22 a_500_n2972# w_n594_n3072# 0.0187f
C23 a_500_n500# w_n594_n600# 0.0187f
C24 a_n500_n3069# a_n500_n4305# 1.03f
C25 w_n594_1872# a_500_736# 0.0023f
C26 a_n500_n597# w_n594_n600# 0.593f
C27 a_n558_1972# a_n558_736# 0.0105f
C28 a_n500_n3069# w_n594_n3072# 0.593f
C29 w_n594_6816# a_n500_6819# 0.593f
C30 a_500_n4208# a_500_n5444# 0.0105f
C31 a_500_n1736# a_n558_n1736# 0.0663f
C32 w_n594_1872# a_n558_736# 0.0023f
C33 a_500_n6680# a_n500_n6777# 0.204f
C34 a_n500_4347# a_n500_3111# 1.03f
C35 w_n594_n4308# a_500_n5444# 0.0023f
C36 a_500_n2972# a_500_n4208# 0.0105f
C37 w_n594_n6780# a_n500_n5541# 0.00575f
C38 a_500_n2972# w_n594_n4308# 0.0023f
C39 a_500_n500# a_n558_n500# 0.0663f
C40 a_n500_n597# a_n558_n500# 0.204f
C41 a_n558_n500# w_n594_n1836# 0.0023f
C42 a_500_n1736# a_n500_n1833# 0.204f
C43 a_500_n6680# a_500_n5444# 0.0105f
C44 a_n558_n4208# a_n558_n5444# 0.0105f
C45 a_n500_n3069# w_n594_n4308# 0.00575f
C46 w_n594_n4308# a_n558_n5444# 0.0023f
C47 w_n594_5580# a_n500_6819# 0.00575f
C48 w_n594_6816# a_n558_6916# 0.0187f
C49 a_n500_8055# a_n558_8152# 0.204f
C50 a_n558_n500# w_n594_636# 0.0023f
C51 w_n594_1872# a_500_3208# 0.0023f
C52 w_n594_3108# a_n558_1972# 0.0023f
C53 w_n594_4344# a_500_5680# 0.0023f
C54 w_n594_5580# a_n500_4347# 0.00575f
C55 w_n594_3108# a_n500_1875# 0.00575f
C56 a_500_n6680# w_n594_n8016# 0.0023f
C57 w_n594_5580# a_n558_6916# 0.0023f
C58 w_n594_4344# a_n558_5680# 0.0023f
C59 a_n558_4444# a_n558_3208# 0.0105f
C60 a_n500_8055# a_n500_6819# 1.03f
C61 a_n558_8152# a_500_8152# 0.0663f
C62 a_n558_n1736# w_n594_n600# 0.0023f
C63 a_n558_n6680# a_500_n6680# 0.0663f
C64 a_500_n9152# a_500_n7916# 0.0105f
C65 a_n500_n4305# w_n594_n5544# 0.00575f
C66 a_500_n9152# a_n558_n9152# 0.0663f
C67 w_n594_5580# a_n558_4444# 0.0023f
C68 a_n500_n9249# w_n594_n9252# 0.593f
C69 a_n500_3111# a_n558_3208# 0.204f
C70 a_n500_n1833# w_n594_n600# 0.00575f
C71 a_n558_n1736# a_n558_n500# 0.0105f
C72 a_n558_n1736# w_n594_n3072# 0.0023f
C73 w_n594_8052# a_n500_8055# 0.593f
C74 a_500_n4208# w_n594_n5544# 0.0023f
C75 a_n558_n4208# w_n594_n5544# 0.0023f
C76 w_n594_4344# a_500_4444# 0.0187f
C77 w_n594_4344# a_n500_5583# 0.00575f
C78 a_500_n1736# w_n594_n600# 0.0023f
C79 a_500_1972# w_n594_636# 0.0023f
C80 a_n558_n2972# w_n594_n3072# 0.0187f
C81 a_n500_n8013# w_n594_n9252# 0.00575f
C82 a_n500_n8013# a_n500_n6777# 1.03f
C83 a_n500_n1833# w_n594_n3072# 0.00575f
C84 a_500_4444# a_500_3208# 0.0105f
C85 w_n594_n8016# a_n500_n6777# 0.00575f
C86 a_500_n6680# w_n594_n5544# 0.0023f
C87 a_n558_1972# a_500_1972# 0.0663f
C88 a_n500_n9249# a_n500_n8013# 1.03f
C89 a_n558_736# a_500_736# 0.0663f
C90 a_500_1972# a_n500_1875# 0.204f
C91 w_n594_8052# a_500_8152# 0.0187f
C92 w_n594_1872# a_500_1972# 0.0187f
C93 a_n500_n9249# w_n594_n8016# 0.00575f
C94 a_n500_n4305# a_n500_n5541# 1.03f
C95 w_n594_3108# a_500_4444# 0.0023f
C96 a_n558_n5444# a_500_n5444# 0.0663f
C97 a_500_n1736# w_n594_n3072# 0.0023f
C98 a_n558_n2972# a_n558_n4208# 0.0105f
C99 a_n558_n6680# a_n500_n6777# 0.204f
C100 a_n500_6819# a_500_6916# 0.204f
C101 a_n558_5680# a_n558_6916# 0.0105f
C102 a_n558_n2972# w_n594_n4308# 0.0023f
C103 a_n500_n3069# a_500_n2972# 0.204f
C104 a_500_736# w_n594_n600# 0.0023f
C105 a_500_n6680# a_500_n7916# 0.0105f
C106 a_500_n6680# w_n594_n6780# 0.0187f
C107 a_n500_639# a_n500_n597# 1.03f
C108 w_n594_6816# a_n500_8055# 0.00575f
C109 a_n558_736# w_n594_n600# 0.0023f
C110 a_n500_1875# a_n500_3111# 1.03f
C111 w_n594_1872# a_n500_3111# 0.00575f
C112 a_n558_4444# a_n558_5680# 0.0105f
C113 w_n594_n4308# a_n500_n5541# 0.00575f
C114 a_n500_639# w_n594_636# 0.593f
C115 a_n500_n8013# w_n594_n8016# 0.593f
C116 a_n500_6819# a_n500_5583# 1.03f
C117 a_n558_6916# a_500_6916# 0.0663f
C118 a_500_n2972# w_n594_n1836# 0.0023f
C119 a_n500_639# a_n500_1875# 1.03f
C120 a_n500_n3069# w_n594_n1836# 0.00575f
C121 a_n558_1972# a_n558_3208# 0.0105f
C122 a_n558_736# a_n558_n500# 0.0105f
C123 w_n594_6816# a_500_8152# 0.0023f
C124 w_n594_8052# a_500_6916# 0.0023f
C125 w_n594_1872# a_n500_639# 0.00575f
C126 a_n558_n6680# a_n558_n5444# 0.0105f
C127 a_n500_4347# a_500_4444# 0.204f
C128 w_n594_1872# a_n558_3208# 0.0023f
C129 a_n558_n6680# w_n594_n8016# 0.0023f
C130 w_n594_n9252# a_n558_n7916# 0.0023f
C131 a_n500_4347# a_n500_5583# 1.03f
C132 w_n594_n5544# a_n500_n6777# 0.00575f
C133 w_n594_4344# a_500_3208# 0.0023f
C134 a_500_n500# a_n500_n597# 0.204f
C135 a_500_n500# w_n594_n1836# 0.0023f
C136 a_n500_n597# w_n594_n1836# 0.00575f
C137 w_n594_6816# a_500_5680# 0.0023f
C138 a_n558_n500# w_n594_n600# 0.0187f
C139 w_n594_6816# a_n558_5680# 0.0023f
C140 a_500_n500# w_n594_636# 0.0023f
C141 a_n558_4444# a_500_4444# 0.0663f
C142 a_n500_n597# w_n594_636# 0.00575f
C143 w_n594_n5544# a_500_n5444# 0.0187f
C144 a_500_n7916# w_n594_n9252# 0.0023f
C145 w_n594_n6780# a_n500_n6777# 0.593f
C146 w_n594_3108# a_500_3208# 0.0187f
C147 a_n558_n9152# w_n594_n9252# 0.0187f
C148 a_n500_n4305# w_n594_n3072# 0.00575f
C149 w_n594_5580# a_500_5680# 0.0187f
C150 a_n500_n9249# a_n558_n9152# 0.204f
C151 a_n500_n8013# a_n558_n7916# 0.204f
C152 w_n594_6816# a_500_6916# 0.0187f
C153 w_n594_n5544# a_n558_n5444# 0.0187f
C154 w_n594_5580# a_n558_5680# 0.0187f
C155 a_n558_1972# w_n594_636# 0.0023f
C156 a_n500_8055# a_500_8152# 0.204f
C157 w_n594_n8016# a_n558_n7916# 0.0187f
C158 a_n500_1875# w_n594_636# 0.00575f
C159 w_n594_n6780# a_500_n5444# 0.0023f
C160 a_n500_n4305# a_500_n4208# 0.204f
C161 a_n500_n4305# a_n558_n4208# 0.204f
C162 a_n500_n4305# w_n594_n4308# 0.593f
C163 a_n500_n5541# a_n500_n6777# 1.03f
C164 a_n558_1972# a_n500_1875# 0.204f
C165 a_500_1972# a_500_736# 0.0105f
C166 w_n594_1872# a_n558_1972# 0.0187f
C167 a_500_n4208# w_n594_n3072# 0.0023f
C168 a_n558_n4208# w_n594_n3072# 0.0023f
C169 w_n594_1872# a_n500_1875# 0.593f
C170 w_n594_4344# a_n500_4347# 0.593f
C171 a_n558_n6680# a_n558_n7916# 0.0105f
C172 a_n558_n6680# w_n594_n5544# 0.0023f
C173 a_n558_n2972# a_500_n2972# 0.0663f
C174 w_n594_6816# a_n500_5583# 0.00575f
C175 w_n594_5580# a_500_6916# 0.0023f
C176 a_500_n7916# a_n500_n8013# 0.204f
C177 w_n594_n6780# a_n558_n5444# 0.0023f
C178 a_n500_n8013# w_n594_n6780# 0.00575f
C179 a_500_n7916# w_n594_n8016# 0.0187f
C180 a_n558_n9152# w_n594_n8016# 0.0023f
C181 a_n500_n3069# a_n558_n2972# 0.204f
C182 a_n500_n5541# a_500_n5444# 0.204f
C183 a_n500_n3069# a_n500_n1833# 1.03f
C184 a_n558_n1736# w_n594_n1836# 0.0187f
C185 a_n558_n4208# a_500_n4208# 0.0663f
C186 a_500_n4208# w_n594_n4308# 0.0187f
C187 a_n558_n4208# w_n594_n4308# 0.0187f
C188 a_500_n1736# a_500_n2972# 0.0105f
C189 w_n594_3108# a_n500_4347# 0.00575f
C190 w_n594_4344# a_n558_4444# 0.0187f
C191 w_n594_5580# a_500_4444# 0.0023f
C192 a_n558_n6680# w_n594_n6780# 0.0187f
C193 w_n594_5580# a_n500_5583# 0.593f
C194 a_n558_8152# a_n558_6916# 0.0105f
C195 a_n500_n5541# a_n558_n5444# 0.204f
C196 a_n558_n2972# w_n594_n1836# 0.0023f
C197 a_n500_n1833# a_n500_n597# 1.03f
C198 a_500_1972# a_500_3208# 0.0105f
C199 a_n500_n1833# w_n594_n1836# 0.593f
C200 a_n500_639# a_500_736# 0.204f
C201 w_n594_8052# a_n558_8152# 0.0187f
C202 w_n594_3108# a_500_1972# 0.0023f
C203 w_n594_4344# a_n500_3111# 0.00575f
C204 w_n594_3108# a_n558_4444# 0.0023f
C205 a_500_n9152# w_n594_n9252# 0.0187f
C206 a_500_n1736# a_500_n500# 0.0105f
C207 a_n500_639# a_n558_736# 0.204f
C208 a_500_5680# a_n558_5680# 0.0663f
C209 a_500_n1736# w_n594_n1836# 0.0187f
C210 a_500_n9152# a_n500_n9249# 0.204f
C211 a_500_8152# a_500_6916# 0.0105f
C212 a_n500_6819# a_n558_6916# 0.204f
C213 a_n500_3111# a_500_3208# 0.204f
C214 w_n594_8052# a_n500_6819# 0.00575f
C215 a_n500_639# w_n594_n600# 0.00575f
C216 a_500_n9152# VSUBS 0.561f
C217 a_n558_n9152# VSUBS 0.561f
C218 a_n500_n9249# VSUBS 1.74f
C219 a_500_n7916# VSUBS 0.548f
C220 a_n558_n7916# VSUBS 0.548f
C221 a_n500_n8013# VSUBS 1.17f
C222 a_500_n6680# VSUBS 0.548f
C223 a_n558_n6680# VSUBS 0.548f
C224 a_n500_n6777# VSUBS 1.17f
C225 a_500_n5444# VSUBS 0.548f
C226 a_n558_n5444# VSUBS 0.548f
C227 a_n500_n5541# VSUBS 1.17f
C228 a_500_n4208# VSUBS 0.548f
C229 a_n558_n4208# VSUBS 0.548f
C230 a_n500_n4305# VSUBS 1.17f
C231 a_500_n2972# VSUBS 0.548f
C232 a_n558_n2972# VSUBS 0.548f
C233 a_n500_n3069# VSUBS 1.17f
C234 a_500_n1736# VSUBS 0.548f
C235 a_n558_n1736# VSUBS 0.548f
C236 a_n500_n1833# VSUBS 1.17f
C237 a_500_n500# VSUBS 0.548f
C238 a_n558_n500# VSUBS 0.548f
C239 a_n500_n597# VSUBS 1.17f
C240 a_500_736# VSUBS 0.548f
C241 a_n558_736# VSUBS 0.548f
C242 a_n500_639# VSUBS 1.17f
C243 a_500_1972# VSUBS 0.548f
C244 a_n558_1972# VSUBS 0.548f
C245 a_n500_1875# VSUBS 1.17f
C246 a_500_3208# VSUBS 0.548f
C247 a_n558_3208# VSUBS 0.548f
C248 a_n500_3111# VSUBS 1.17f
C249 a_500_4444# VSUBS 0.548f
C250 a_n558_4444# VSUBS 0.548f
C251 a_n500_4347# VSUBS 1.17f
C252 a_500_5680# VSUBS 0.548f
C253 a_n558_5680# VSUBS 0.548f
C254 a_n500_5583# VSUBS 1.17f
C255 a_500_6916# VSUBS 0.548f
C256 a_n558_6916# VSUBS 0.548f
C257 a_n500_6819# VSUBS 1.17f
C258 a_500_8152# VSUBS 0.561f
C259 a_n558_8152# VSUBS 0.561f
C260 a_n500_8055# VSUBS 1.74f
C261 w_n594_n9252# VSUBS 4.28f
C262 w_n594_n8016# VSUBS 4.28f
C263 w_n594_n6780# VSUBS 4.28f
C264 w_n594_n5544# VSUBS 4.28f
C265 w_n594_n4308# VSUBS 4.28f
C266 w_n594_n3072# VSUBS 4.28f
C267 w_n594_n1836# VSUBS 4.28f
C268 w_n594_n600# VSUBS 4.28f
C269 w_n594_636# VSUBS 4.28f
C270 w_n594_1872# VSUBS 4.28f
C271 w_n594_3108# VSUBS 4.28f
C272 w_n594_4344# VSUBS 4.28f
C273 w_n594_5580# VSUBS 4.28f
C274 w_n594_6816# VSUBS 4.28f
C275 w_n594_8052# VSUBS 4.28f
.ends

.subckt sky130_fd_pr__nfet_01v8_3ZAA45 a_100_n500# a_n158_n500# a_n100_n588# VSUBS
X0 a_100_n500# a_n100_n588# a_n158_n500# VSUBS sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=1
**devattr s=58000,2116 d=58000,2116
C0 a_n100_n588# a_100_n500# 0.112f
C1 a_n100_n588# a_n158_n500# 0.112f
C2 a_n158_n500# a_100_n500# 0.274f
C3 a_100_n500# VSUBS 0.505f
C4 a_n158_n500# VSUBS 0.505f
C5 a_n100_n588# VSUBS 0.687f
.ends

.subckt sky130_fd_pr__pfet_01v8_SKU9VM a_n500_n597# a_500_n500# w_n594_n600# a_n558_n500#
+ VSUBS
X0 a_500_n500# a_n500_n597# a_n558_n500# w_n594_n600# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
C0 w_n594_n600# a_n558_n500# 0.0187f
C1 a_500_n500# w_n594_n600# 0.0187f
C2 a_500_n500# a_n558_n500# 0.0663f
C3 w_n594_n600# a_n500_n597# 0.593f
C4 a_n500_n597# a_n558_n500# 0.204f
C5 a_500_n500# a_n500_n597# 0.204f
C6 a_500_n500# VSUBS 0.573f
C7 a_n558_n500# VSUBS 0.573f
C8 a_n500_n597# VSUBS 2.31f
C9 w_n594_n600# VSUBS 4.28f
.ends

.subckt sky130_fd_pr__pfet_01v8_E769TZ a_n1558_11242# a_n1558_n14714# a_n1500_n43239#
+ w_n1594_n3690# a_n1500_n11103# a_n1558_50794# a_1500_n23366# a_n1500_n50655# w_n1594_n56838#
+ w_n1594_n24702# a_1500_n30782# a_n1500_3729# a_n1558_n60446# w_n1594_12378# w_n1594_n63018#
+ a_1500_n8534# a_n1558_14950# a_1500_n19658# a_n1500_n14811# a_n1500_n46947# w_n1594_9906#
+ w_n1594_n6162# a_1500_22366# a_n1500_22269# a_n1558_53266# a_n1558_n56738# a_n1558_n24602#
+ a_n1558_21130# a_n1500_n53127# w_n1594_n13578# a_n1558_60682# a_1500_n33254# a_n1500_n60543#
+ w_n1594_n20994# a_1500_n40670# a_1500_18658# a_n1558_49558# a_n1558_17422# w_n1594_22266#
+ a_n1500_n49419# w_n1594_n9870# a_n1500_25977# a_n1558_56974# a_n1500_n56835# a_1500_n29546#
+ a_n1558_n3590# a_1500_n36962# a_n1500_9909# a_n1558_n13478# a_1500_32254# a_n1500_32157#
+ a_n1558_n20894# a_n1500_n63015# w_n1594_18558# w_n1594_n23466# a_1500_n43142# w_n1594_n30882#
+ w_n1594_25974# a_n1500_n2451# a_1500_28546# a_1500_n7298# a_n1500_28449# a_n1558_59446#
+ a_n1558_27310# a_n1500_n13575# a_n1500_n59307# w_n1594_32154# w_n1594_n19758# a_1500_35962#
+ a_n1558_n6062# a_n1500_35865# a_1500_n39434# a_n1500_n20991# a_n1558_n23366# a_1500_n46850#
+ a_1500_42142# a_n1500_42045# a_n1558_n30782# w_n1594_n33354# w_n1594_28446# a_1500_n53030#
+ w_n1594_n40770# w_n1594_35862# a_n1558_n9770# w_n1594_18# a_n1558_16186# a_n1500_21#
+ a_n1558_n19658# a_n1500_n16047# a_1500_38434# a_n1500_38337# a_n1500_n55599# a_n1500_n23463#
+ w_n1594_n29646# a_1500_45850# w_n1594_42042# a_n1500_45753# a_n1558_40906# a_1500_n49322#
+ a_n1558_n33254# a_1500_52030# a_n1500_n8631# a_n1558_n40670# a_n1558_19894# w_n1594_n43242#
+ a_n1500_n19755# w_n1594_38334# w_n1594_45750# a_n1558_26074# a_n1558_n29546# a_1500_48322#
+ a_n1500_48225# a_1500_n38198# a_n1558_33490# a_n1558_n36962# a_n1500_n33351# w_n1594_n39534#
+ a_n1500_55641# a_1500_n59210# w_n1594_n46950# a_1500_n62918# a_n1558_n43142# a_n1558_29782#
+ w_n1594_n53130# a_n1500_n29643# w_n1594_48222# a_1500_37198# a_n1558_n39434# a_1500_58210#
+ a_n1500_58113# a_n1500_12381# a_1500_n1118# a_1500_n48086# a_n1558_n46850# a_1500_61918#
+ w_n1594_n49422# a_n1500_n7395# a_n1558_n53030# w_n1594_37098# a_n1558_39670# a_n1500_n39531#
+ w_n1594_58110# a_1500_n4826# w_n1594_61818# a_1500_47086# a_n1558_10006# a_n1558_n49322#
+ w_n1594_n2454# w_n1594_n38298# a_1500_2590# w_n1594_2490# w_n1594_n59310# a_n1500_6201#
+ a_n1500_18561# a_n1558_13714# a_n1558_2590# a_1500_n25838# a_n1558_n38198# a_1500_5062#
+ a_1500_118# a_n1558_n59210# w_n1594_n48186# w_n1594_n16050# a_n1558_n62918# a_1500_n32018#
+ a_n1500_2493# a_1500_24838# a_n1558_5062# a_n1500_n38295# w_n1594_n8634# a_1500_8770#
+ a_n1558_55738# a_n1558_23602# a_n1558_n2354# w_n1594_8670# a_1500_n35726# a_n1558_n48086#
+ a_1500_31018# w_n1594_n58074# w_n1594_24738# a_n1558_8770# a_n1500_n1215# a_n1558_12478#
+ a_n1500_n12339# a_n1500_n48183# a_1500_34726# a_n1500_34629# w_n1594_n25938# a_1500_n45614#
+ a_n1500_8673# w_n1594_n32118# a_n1500_n4923# w_n1594_34626# a_n1558_n8534# w_n1594_n7398#
+ a_n1558_22366# a_n1558_n25838# a_n1500_n22227# a_n1500_n58071# a_1500_44614# a_n1500_44517#
+ a_n1500_n61779# w_n1594_n35826# a_n1500_51933# a_1500_n55502# a_n1558_n32018# a_n1558_18658#
+ w_n1594_n42006# a_n1500_n18519# a_n1500_n25935# w_n1594_44514# w_n1594_51930# a_n1558_32254#
+ a_n1558_n35726# a_n1500_n32115# a_1500_54502# a_n1500_54405# a_1500_n44378# a_1500_n12242#
+ w_n1594_n45714# a_n1500_61821# a_1500_n51794# a_n1500_n3687# a_n1558_28546# a_n1558_n7298#
+ a_n1500_n28407# a_n1558_35962# a_n1500_n35823# w_n1594_54402# a_1500_n15950# a_1500_43378#
+ a_1500_11242# a_n1500_11145# a_n1558_42142# a_n1558_n45614# a_1500_50794# a_n1500_n42003#
+ a_n1500_50697# a_1500_n54266# a_1500_n22130# a_n1500_n6159# w_n1594_n55602# a_1500_n61682#
+ a_n1558_38434# a_n1500_n24699# w_n1594_43278# w_n1594_11142# a_1500_14950# a_n1500_46989#
+ a_n1558_45850# a_n1500_14853# a_1500_n18422# a_n1500_n45711# w_n1594_50694# a_1500_n57974#
+ a_n1500_n9867# w_n1594_n1218# a_1500_53266# a_1500_1354# a_n1500_53169# a_1500_21130#
+ a_n1500_21033# a_n1558_n55502# a_n1558_52030# w_n1594_1254# w_n1594_n12342# w_n1594_n44478#
+ a_1500_60682# a_n1500_60585# w_n1594_14850# w_n1594_n51894# w_n1594_46986# a_1500_49558#
+ a_1500_17422# a_n1558_48322# a_n1500_17325# a_n1500_n34587# a_1500_56974# a_n1558_1354#
+ w_n1594_53166# w_n1594_21030# w_n1594_n4926# a_n1500_56877# a_n1500_24741# a_1500_n3590#
+ a_1500_n28310# w_n1594_60582# w_n1594_4962# a_n1558_n44378# a_n1558_n12242# a_n1558_n51794#
+ w_n1594_17322# w_n1594_n22230# w_n1594_n54366# w_n1594_49458# a_n1500_1257# w_n1594_n61782#
+ w_n1594_56874# a_n1558_37198# a_n1500_n37059# a_1500_59446# a_1500_27310# a_1500_7534#
+ a_n1500_59349# a_n1500_27213# a_1500_n6062# a_1500_n17186# a_n1558_58210# a_n1558_n15950#
+ a_n1500_n44475# a_n1558_n1118# w_n1594_7434# w_n1594_n18522# a_n1558_61918# a_n1500_n51891#
+ a_n1558_n54266# a_1500_n41906# a_n1500_4965# a_n1558_n22130# a_n1558_n61682# w_n1594_59346#
+ w_n1594_27210# a_n1558_7534# a_1500_n9770# w_n1594_30918# a_n1558_n4826# a_1500_16186#
+ a_n1500_16089# a_n1558_47086# a_n1558_n18422# a_n1500_37101# a_n1558_n57974# a_1500_n27074#
+ a_n1500_n54363# a_1500_40906# w_n1594_n28410# a_n1500_40809# a_1500_n34490# a_n1500_7437#
+ w_n1594_16086# a_1500_19894# a_n1500_19797# w_n1594_40806# a_1500_26074# a_1500_6298#
+ a_n1558_n28310# w_n1594_6198# w_n1594_n17286# a_1500_33490# a_n1500_33393# w_n1594_19794#
+ a_n1558_6298# a_1500_29782# a_n1500_29685# a_n1558_24838# w_n1594_33390# a_n1558_n17186#
+ a_n1558_118# a_n1558_31018# w_n1594_n27174# a_n1500_43281# a_n1558_n41906# a_1500_n11006#
+ w_n1594_29682# w_n1594_n34590# a_1500_n50558# a_n1500_n17283# a_1500_39670# a_n1500_39573#
+ a_n1558_34726# a_1500_n14714# a_n1558_n27074# a_1500_10006# a_n1558_n34490# w_n1594_n37062#
+ w_n1594_39570# a_1500_n60446# a_n1500_n27171# a_1500_13714# a_n1500_13617# a_n1500_49461#
+ a_n1558_44614# a_n1500_n30879# a_1500_n56738# a_1500_n24602# w_n1594_n11106# w_n1594_n50658#
+ w_n1594_13614# a_1500_55738# a_1500_23602# a_1500_3826# a_n1500_23505# a_1500_n2354#
+ a_1500_n13478# a_n1558_54502# a_n1500_n40767# w_n1594_3726# w_n1594_n14814# a_n1500_30921#
+ a_1500_n20894# a_n1558_n11006# a_n1558_n50558# w_n1594_n60546# a_n1558_3826# w_n1594_55638#
+ w_n1594_23502# VSUBS a_1500_12478# a_n1558_43378#
X0 a_1500_53266# a_n1500_53169# a_n1558_53266# w_n1594_53166# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X1 a_1500_n18422# a_n1500_n18519# a_n1558_n18422# w_n1594_n18522# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X2 a_1500_n45614# a_n1500_n45711# a_n1558_n45614# w_n1594_n45714# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X3 a_1500_n43142# a_n1500_n43239# a_n1558_n43142# w_n1594_n43242# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X4 a_1500_n22130# a_n1500_n22227# a_n1558_n22130# w_n1594_n22230# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X5 a_1500_n3590# a_n1500_n3687# a_n1558_n3590# w_n1594_n3690# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X6 a_1500_35962# a_n1500_35865# a_n1558_35962# w_n1594_35862# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X7 a_1500_33490# a_n1500_33393# a_n1558_33490# w_n1594_33390# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X8 a_1500_60682# a_n1500_60585# a_n1558_60682# w_n1594_60582# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X9 a_1500_12478# a_n1500_12381# a_n1558_12478# w_n1594_12378# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X10 a_1500_38434# a_n1500_38337# a_n1558_38434# w_n1594_38334# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X11 a_1500_6298# a_n1500_6201# a_n1558_6298# w_n1594_6198# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X12 a_1500_n55502# a_n1500_n55599# a_n1558_n55502# w_n1594_n55602# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X13 a_1500_n32018# a_n1500_n32115# a_n1558_n32018# w_n1594_n32118# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X14 a_1500_45850# a_n1500_45753# a_n1558_45850# w_n1594_45750# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X15 a_1500_24838# a_n1500_24741# a_n1558_24838# w_n1594_24738# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X16 a_1500_n38198# a_n1500_n38295# a_n1558_n38198# w_n1594_n38298# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X17 a_1500_22366# a_n1500_22269# a_n1558_22366# w_n1594_22266# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X18 a_1500_48322# a_n1500_48225# a_n1558_48322# w_n1594_48222# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X19 a_1500_n14714# a_n1500_n14811# a_n1558_n14714# w_n1594_n14814# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X20 a_1500_n41906# a_n1500_n42003# a_n1558_n41906# w_n1594_n42006# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X21 a_1500_n12242# a_n1500_n12339# a_n1558_n12242# w_n1594_n12342# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X22 a_1500_34726# a_n1500_34629# a_n1558_34726# w_n1594_34626# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X23 a_1500_61918# a_n1500_61821# a_n1558_61918# w_n1594_61818# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X24 a_1500_32254# a_n1500_32157# a_n1558_32254# w_n1594_32154# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X25 a_1500_n48086# a_n1500_n48183# a_n1558_n48086# w_n1594_n48186# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X26 a_1500_58210# a_n1500_58113# a_n1558_58210# w_n1594_58110# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X27 a_1500_n24602# a_n1500_n24699# a_n1558_n24602# w_n1594_n24702# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X28 a_1500_14950# a_n1500_14853# a_n1558_14950# w_n1594_14850# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X29 a_1500_n8534# a_n1500_n8631# a_n1558_n8534# w_n1594_n8634# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X30 a_1500_n57974# a_n1500_n58071# a_n1558_n57974# w_n1594_n58074# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X31 a_1500_n6062# a_n1500_n6159# a_n1558_n6062# w_n1594_n6162# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X32 a_1500_n34490# a_n1500_n34587# a_n1558_n34490# w_n1594_n34590# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X33 a_1500_17422# a_n1500_17325# a_n1558_17422# w_n1594_17322# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X34 a_1500_44614# a_n1500_44517# a_n1558_44614# w_n1594_44514# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X35 a_1500_42142# a_n1500_42045# a_n1558_42142# w_n1594_42042# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X36 a_1500_8770# a_n1500_8673# a_n1558_8770# w_n1594_8670# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X37 a_1500_n11006# a_n1500_n11103# a_n1558_n11006# w_n1594_n11106# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X38 a_1500_n19658# a_n1500_n19755# a_n1558_n19658# w_n1594_n19758# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X39 a_1500_n46850# a_n1500_n46947# a_n1558_n46850# w_n1594_n46950# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X40 a_1500_n17186# a_n1500_n17283# a_n1558_n17186# w_n1594_n17286# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X41 a_1500_27310# a_n1500_27213# a_n1558_27310# w_n1594_27210# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X42 a_1500_n44378# a_n1500_n44475# a_n1558_n44378# w_n1594_n44478# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X43 a_1500_54502# a_n1500_54405# a_n1558_54502# w_n1594_54402# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X44 a_1500_52030# a_n1500_51933# a_n1558_52030# w_n1594_51930# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X45 a_1500_31018# a_n1500_30921# a_n1558_31018# w_n1594_30918# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X46 a_1500_n4826# a_n1500_n4923# a_n1558_n4826# w_n1594_n4926# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X47 a_1500_37198# a_n1500_37101# a_n1558_37198# w_n1594_37098# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X48 a_1500_n2354# a_n1500_n2451# a_n1558_n2354# w_n1594_n2454# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X49 a_1500_n51794# a_n1500_n51891# a_n1558_n51794# w_n1594_n51894# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X50 a_1500_n29546# a_n1500_n29643# a_n1558_n29546# w_n1594_n29646# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X51 a_1500_13714# a_n1500_13617# a_n1558_13714# w_n1594_13614# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X52 a_1500_n56738# a_n1500_n56835# a_n1558_n56738# w_n1594_n56838# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X53 a_1500_11242# a_n1500_11145# a_n1558_11242# w_n1594_11142# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X54 a_1500_40906# a_n1500_40809# a_n1558_40906# w_n1594_40806# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X55 a_1500_n27074# a_n1500_n27171# a_n1558_n27074# w_n1594_n27174# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X56 a_1500_n54266# a_n1500_n54363# a_n1558_n54266# w_n1594_n54366# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X57 a_1500_19894# a_n1500_19797# a_n1558_19894# w_n1594_19794# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X58 a_1500_2590# a_n1500_2493# a_n1558_2590# w_n1594_2490# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X59 a_1500_n59210# a_n1500_n59307# a_n1558_n59210# w_n1594_n59310# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X60 a_1500_7534# a_n1500_7437# a_n1558_7534# w_n1594_7434# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X61 a_1500_49558# a_n1500_49461# a_n1558_49558# w_n1594_49458# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X62 a_1500_n36962# a_n1500_n37059# a_n1558_n36962# w_n1594_n37062# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X63 a_1500_5062# a_n1500_4965# a_n1558_5062# w_n1594_4962# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X64 a_1500_47086# a_n1500_46989# a_n1558_47086# w_n1594_46986# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X65 a_1500_n15950# a_n1500_n16047# a_n1558_n15950# w_n1594_n16050# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X66 a_1500_n61682# a_n1500_n61779# a_n1558_n61682# w_n1594_n61782# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X67 a_1500_n13478# a_n1500_n13575# a_n1558_n13478# w_n1594_n13578# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X68 a_1500_23602# a_n1500_23505# a_n1558_23602# w_n1594_23502# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X69 a_1500_n40670# a_n1500_n40767# a_n1558_n40670# w_n1594_n40770# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X70 a_1500_n39434# a_n1500_n39531# a_n1558_n39434# w_n1594_n39534# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X71 a_1500_21130# a_n1500_21033# a_n1558_21130# w_n1594_21030# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X72 a_1500_29782# a_n1500_29685# a_n1558_29782# w_n1594_29682# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X73 a_1500_56974# a_n1500_56877# a_n1558_56974# w_n1594_56874# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X74 a_1500_59446# a_n1500_59349# a_n1558_59446# w_n1594_59346# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X75 a_1500_n20894# a_n1500_n20991# a_n1558_n20894# w_n1594_n20994# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X76 a_1500_n25838# a_n1500_n25935# a_n1558_n25838# w_n1594_n25938# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X77 a_1500_n23366# a_n1500_n23463# a_n1558_n23366# w_n1594_n23466# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X78 a_1500_n50558# a_n1500_n50655# a_n1558_n50558# w_n1594_n50658# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X79 a_1500_n49322# a_n1500_n49419# a_n1558_n49322# w_n1594_n49422# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X80 a_1500_n1118# a_n1500_n1215# a_n1558_n1118# w_n1594_n1218# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X81 a_1500_n9770# a_n1500_n9867# a_n1558_n9770# w_n1594_n9870# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X82 a_1500_n28310# a_n1500_n28407# a_n1558_n28310# w_n1594_n28410# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X83 a_1500_n7298# a_n1500_n7395# a_n1558_n7298# w_n1594_n7398# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X84 a_1500_10006# a_n1500_9909# a_n1558_10006# w_n1594_9906# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X85 a_1500_39670# a_n1500_39573# a_n1558_39670# w_n1594_39570# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X86 a_1500_18658# a_n1500_18561# a_n1558_18658# w_n1594_18558# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X87 a_1500_n53030# a_n1500_n53127# a_n1558_n53030# w_n1594_n53130# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X88 a_1500_3826# a_n1500_3729# a_n1558_3826# w_n1594_3726# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X89 a_1500_16186# a_n1500_16089# a_n1558_16186# w_n1594_16086# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X90 a_1500_1354# a_n1500_1257# a_n1558_1354# w_n1594_1254# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X91 a_1500_43378# a_n1500_43281# a_n1558_43378# w_n1594_43278# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X92 a_1500_n30782# a_n1500_n30879# a_n1558_n30782# w_n1594_n30882# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X93 a_1500_118# a_n1500_21# a_n1558_118# w_n1594_18# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X94 a_1500_n35726# a_n1500_n35823# a_n1558_n35726# w_n1594_n35826# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X95 a_1500_n62918# a_n1500_n63015# a_n1558_n62918# w_n1594_n63018# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X96 a_1500_n33254# a_n1500_n33351# a_n1558_n33254# w_n1594_n33354# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X97 a_1500_n60446# a_n1500_n60543# a_n1558_n60446# w_n1594_n60546# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X98 a_1500_50794# a_n1500_50697# a_n1558_50794# w_n1594_50694# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X99 a_1500_28546# a_n1500_28449# a_n1558_28546# w_n1594_28446# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X100 a_1500_55738# a_n1500_55641# a_n1558_55738# w_n1594_55638# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
X101 a_1500_26074# a_n1500_25977# a_n1558_26074# w_n1594_25974# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
C0 w_n1594_54402# a_n1500_55641# 0.0172f
C1 a_n1500_n63015# a_n1558_n62918# 0.217f
C2 w_n1594_17322# a_n1558_16186# 0.0023f
C3 a_1500_n61682# a_1500_n62918# 0.0105f
C4 w_n1594_61818# a_1500_61918# 0.0187f
C5 a_n1500_n45711# w_n1594_n44478# 0.0172f
C6 a_n1500_n28407# a_n1500_n27171# 3.11f
C7 w_n1594_n18522# a_n1558_n19658# 0.0023f
C8 w_n1594_49458# a_n1500_48225# 0.0172f
C9 w_n1594_2490# a_n1500_3729# 0.0172f
C10 a_1500_8770# w_n1594_8670# 0.0187f
C11 w_n1594_55638# a_n1500_55641# 1.65f
C12 w_n1594_n58074# a_n1500_n56835# 0.0172f
C13 w_n1594_n60546# a_1500_n61682# 0.0023f
C14 a_1500_n15950# a_1500_n14714# 0.0105f
C15 a_n1558_6298# w_n1594_7434# 0.0023f
C16 w_n1594_n38298# a_n1558_n36962# 0.0023f
C17 w_n1594_n18522# a_n1558_n17186# 0.0023f
C18 a_n1558_n55502# w_n1594_n56838# 0.0023f
C19 a_n1558_n18422# w_n1594_n17286# 0.0023f
C20 w_n1594_n19758# a_n1500_n20991# 0.0172f
C21 a_n1558_n8534# a_n1558_n7298# 0.0105f
C22 a_1500_n2354# w_n1594_n1218# 0.0023f
C23 w_n1594_n34590# a_1500_n35726# 0.0023f
C24 a_n1500_n30879# w_n1594_n32118# 0.0172f
C25 a_n1500_4965# a_n1500_3729# 3.11f
C26 a_n1500_n30879# w_n1594_n30882# 1.65f
C27 w_n1594_n19758# a_1500_n20894# 0.0023f
C28 a_1500_n6062# a_1500_n7298# 0.0105f
C29 a_n1558_n7298# w_n1594_n7398# 0.0187f
C30 w_n1594_n12342# a_n1500_n12339# 1.65f
C31 a_1500_n23366# a_1500_n24602# 0.0105f
C32 a_n1500_n24699# a_n1558_n24602# 0.217f
C33 a_1500_17422# a_1500_16186# 0.0105f
C34 a_1500_59446# a_1500_60682# 0.0105f
C35 w_n1594_n43242# a_n1558_n44378# 0.0023f
C36 w_n1594_48222# a_n1500_46989# 0.0172f
C37 a_1500_n1118# a_n1500_n1215# 0.217f
C38 a_n1558_24838# a_n1558_26074# 0.0105f
C39 w_n1594_3726# a_1500_2590# 0.0023f
C40 a_n1500_n4923# a_n1500_n6159# 3.11f
C41 w_n1594_n40770# a_n1558_n39434# 0.0023f
C42 w_n1594_16086# a_n1558_17422# 0.0023f
C43 a_1500_19894# w_n1594_19794# 0.0187f
C44 a_n1500_22269# a_n1558_22366# 0.217f
C45 w_n1594_1254# a_n1558_118# 0.0023f
C46 w_n1594_n59310# a_n1500_n58071# 0.0172f
C47 a_n1558_37198# w_n1594_37098# 0.0187f
C48 a_n1500_n4923# w_n1594_n3690# 0.0172f
C49 a_n1500_n48183# a_n1558_n48086# 0.217f
C50 a_n1500_n13575# a_n1558_n13478# 0.217f
C51 a_1500_n46850# a_1500_n48086# 0.0105f
C52 a_n1500_n49419# w_n1594_n50658# 0.0172f
C53 w_n1594_9906# a_n1500_11145# 0.0172f
C54 w_n1594_n4926# a_n1500_n3687# 0.0172f
C55 a_n1558_40906# a_n1500_40809# 0.217f
C56 w_n1594_n38298# a_n1558_n39434# 0.0023f
C57 a_n1500_29685# a_n1500_30921# 3.11f
C58 a_n1500_50697# w_n1594_51930# 0.0172f
C59 w_n1594_n44478# a_n1500_n44475# 1.65f
C60 a_n1500_58113# w_n1594_58110# 1.65f
C61 a_n1500_7437# w_n1594_6198# 0.0172f
C62 w_n1594_55638# a_n1558_56974# 0.0023f
C63 a_n1558_n29546# w_n1594_n28410# 0.0023f
C64 a_1500_33490# w_n1594_34626# 0.0023f
C65 a_n1500_35865# a_n1558_35962# 0.217f
C66 w_n1594_n13578# a_n1500_n13575# 1.65f
C67 a_n1500_22269# a_1500_22366# 0.217f
C68 a_n1558_n44378# a_n1558_n43142# 0.0105f
C69 a_n1500_54405# w_n1594_53166# 0.0172f
C70 a_n1558_37198# w_n1594_35862# 0.0023f
C71 w_n1594_50694# a_n1500_49461# 0.0172f
C72 a_n1558_n57974# a_n1558_n59210# 0.0105f
C73 w_n1594_60582# a_1500_59446# 0.0023f
C74 a_n1558_8770# a_n1558_7534# 0.0105f
C75 a_n1558_39670# a_n1558_38434# 0.0105f
C76 a_n1500_1257# a_n1500_21# 3.11f
C77 w_n1594_n43242# a_n1558_n43142# 0.0187f
C78 a_n1558_10006# a_n1500_9909# 0.217f
C79 w_n1594_n61782# a_1500_n60446# 0.0023f
C80 a_n1558_39670# w_n1594_40806# 0.0023f
C81 a_n1500_58113# a_n1558_58210# 0.217f
C82 a_n1558_n54266# a_n1558_n55502# 0.0105f
C83 a_1500_n6062# w_n1594_n7398# 0.0023f
C84 a_1500_n11006# a_n1500_n11103# 0.217f
C85 a_1500_8770# w_n1594_7434# 0.0023f
C86 w_n1594_n55602# a_n1558_n56738# 0.0023f
C87 w_n1594_17322# a_n1500_16089# 0.0172f
C88 w_n1594_n25938# a_n1558_n25838# 0.0187f
C89 w_n1594_16086# a_1500_17422# 0.0023f
C90 a_n1558_n45614# w_n1594_n45714# 0.0187f
C91 a_n1558_n25838# w_n1594_n24702# 0.0023f
C92 a_1500_n11006# w_n1594_n11106# 0.0187f
C93 a_n1558_n50558# w_n1594_n49422# 0.0023f
C94 w_n1594_60582# a_n1558_59446# 0.0023f
C95 a_n1558_40906# w_n1594_42042# 0.0023f
C96 a_n1500_34629# a_1500_34726# 0.217f
C97 a_n1500_n39531# a_n1500_n40767# 3.11f
C98 a_n1500_17325# a_n1558_17422# 0.217f
C99 a_n1500_n7395# w_n1594_n6162# 0.0172f
C100 a_n1500_n2451# w_n1594_n3690# 0.0172f
C101 w_n1594_19794# a_n1500_19797# 1.65f
C102 a_n1500_6201# a_1500_6298# 0.217f
C103 a_n1558_n55502# w_n1594_n54366# 0.0023f
C104 w_n1594_n56838# a_n1558_n57974# 0.0023f
C105 w_n1594_n60546# a_1500_n60446# 0.0187f
C106 a_1500_19894# w_n1594_18558# 0.0023f
C107 w_n1594_n29646# a_1500_n28310# 0.0023f
C108 a_n1500_n33351# a_n1558_n33254# 0.217f
C109 a_n1500_n3687# w_n1594_n3690# 1.65f
C110 w_n1594_4962# a_n1558_5062# 0.0187f
C111 a_n1500_55641# a_1500_55738# 0.217f
C112 w_n1594_n34590# a_1500_n34490# 0.0187f
C113 a_n1500_n20991# a_1500_n20894# 0.217f
C114 a_1500_50794# a_1500_52030# 0.0105f
C115 w_n1594_n33354# a_1500_n34490# 0.0023f
C116 a_n1500_n43239# a_1500_n43142# 0.217f
C117 a_n1500_n29643# w_n1594_n30882# 0.0172f
C118 w_n1594_61818# a_n1500_60585# 0.0172f
C119 w_n1594_50694# a_n1500_51933# 0.0172f
C120 a_n1500_n29643# a_n1500_n28407# 3.11f
C121 w_n1594_18# a_n1558_n1118# 0.0023f
C122 a_n1500_56877# w_n1594_55638# 0.0172f
C123 a_n1558_6298# w_n1594_6198# 0.0187f
C124 a_n1500_30921# a_n1558_31018# 0.217f
C125 w_n1594_33390# a_n1500_32157# 0.0172f
C126 a_n1500_1257# a_1500_1354# 0.217f
C127 a_n1500_42045# a_n1500_40809# 3.11f
C128 w_n1594_59346# a_n1500_60585# 0.0172f
C129 w_n1594_n38298# a_n1558_n38198# 0.0187f
C130 a_1500_32254# w_n1594_30918# 0.0023f
C131 w_n1594_n13578# a_n1500_n12339# 0.0172f
C132 w_n1594_45750# a_1500_45850# 0.0187f
C133 w_n1594_40806# a_n1500_40809# 1.65f
C134 w_n1594_n44478# a_n1500_n43239# 0.0172f
C135 a_1500_32254# a_n1500_32157# 0.217f
C136 w_n1594_9906# a_n1500_8673# 0.0172f
C137 w_n1594_1254# a_1500_2590# 0.0023f
C138 a_1500_17422# a_n1500_17325# 0.217f
C139 a_n1558_n11006# w_n1594_n9870# 0.0023f
C140 a_n1500_n50655# a_n1500_n51891# 3.11f
C141 a_n1500_n8631# a_n1500_n9867# 3.11f
C142 a_n1500_34629# w_n1594_35862# 0.0172f
C143 a_n1500_n6159# w_n1594_n6162# 1.65f
C144 a_n1500_23505# w_n1594_22266# 0.0172f
C145 w_n1594_n13578# a_1500_n14714# 0.0023f
C146 a_n1500_n2451# a_n1500_n1215# 3.11f
C147 a_n1558_27310# w_n1594_25974# 0.0023f
C148 a_n1500_25977# w_n1594_27210# 0.0172f
C149 w_n1594_2490# a_1500_3826# 0.0023f
C150 a_n1558_22366# w_n1594_23502# 0.0023f
C151 w_n1594_n4926# a_1500_n3590# 0.0023f
C152 a_n1500_n58071# a_1500_n57974# 0.217f
C153 a_n1558_n24602# w_n1594_n25938# 0.0023f
C154 a_n1558_n4826# a_n1558_n6062# 0.0105f
C155 a_n1558_n24602# w_n1594_n24702# 0.0187f
C156 w_n1594_9906# a_n1500_9909# 1.65f
C157 a_n1558_n55502# a_n1558_n56738# 0.0105f
C158 w_n1594_19794# a_n1558_19894# 0.0187f
C159 w_n1594_n42006# a_n1558_n43142# 0.0023f
C160 w_n1594_n43242# a_n1558_n41906# 0.0023f
C161 a_n1558_28546# w_n1594_27210# 0.0023f
C162 a_n1500_n54363# a_1500_n54266# 0.217f
C163 a_n1558_21130# w_n1594_19794# 0.0023f
C164 w_n1594_18558# a_n1500_19797# 0.0172f
C165 a_1500_28546# w_n1594_27210# 0.0023f
C166 a_n1558_n44378# w_n1594_n45714# 0.0023f
C167 w_n1594_n37062# a_1500_n35726# 0.0023f
C168 a_n1558_3826# a_n1558_5062# 0.0105f
C169 w_n1594_50694# a_n1558_52030# 0.0023f
C170 a_n1558_n49322# w_n1594_n49422# 0.0187f
C171 a_n1500_42045# w_n1594_42042# 1.65f
C172 w_n1594_32154# a_1500_32254# 0.0187f
C173 a_n1500_n61779# a_n1558_n61682# 0.217f
C174 a_1500_n60446# a_1500_n61682# 0.0105f
C175 w_n1594_n19758# a_n1500_n18519# 0.0172f
C176 a_n1558_n54266# w_n1594_n53130# 0.0023f
C177 w_n1594_60582# a_n1558_61918# 0.0023f
C178 w_n1594_58110# a_n1500_59349# 0.0172f
C179 a_1500_22366# w_n1594_23502# 0.0023f
C180 a_1500_19894# a_1500_21130# 0.0105f
C181 a_n1500_58113# a_1500_58210# 0.217f
C182 w_n1594_n60546# a_1500_n59210# 0.0023f
C183 a_n1558_n54266# w_n1594_n54366# 0.0187f
C184 w_n1594_n56838# a_n1558_n56738# 0.0187f
C185 a_n1558_44614# w_n1594_44514# 0.0187f
C186 a_1500_n48086# w_n1594_n46950# 0.0023f
C187 w_n1594_n34590# a_1500_n33254# 0.0023f
C188 a_n1500_12381# a_n1500_13617# 3.11f
C189 w_n1594_50694# a_1500_52030# 0.0023f
C190 w_n1594_n33354# a_1500_n33254# 0.0187f
C191 a_1500_54502# a_n1500_54405# 0.217f
C192 a_n1500_39573# w_n1594_40806# 0.0172f
C193 a_n1558_n41906# a_n1558_n43142# 0.0105f
C194 w_n1594_n37062# a_1500_n38198# 0.0023f
C195 w_n1594_n35826# a_1500_n35726# 0.0187f
C196 a_n1558_1354# w_n1594_2490# 0.0023f
C197 w_n1594_12378# a_1500_11242# 0.0023f
C198 w_n1594_8670# a_n1500_8673# 1.65f
C199 a_1500_n7298# w_n1594_n6162# 0.0023f
C200 a_n1500_n30879# a_n1500_n32115# 3.11f
C201 w_n1594_58110# a_n1558_56974# 0.0023f
C202 w_n1594_n32118# a_n1500_n33351# 0.0172f
C203 w_n1594_24738# a_1500_26074# 0.0023f
C204 a_1500_3826# a_1500_5062# 0.0105f
C205 a_n1500_14853# a_n1558_14950# 0.217f
C206 a_n1500_n9867# w_n1594_n9870# 1.65f
C207 a_n1500_n35823# a_n1500_n37059# 3.11f
C208 a_1500_n49322# w_n1594_n48186# 0.0023f
C209 a_1500_n45614# a_1500_n46850# 0.0105f
C210 a_n1500_n46947# a_n1558_n46850# 0.217f
C211 w_n1594_n27174# a_n1558_n28310# 0.0023f
C212 w_n1594_12378# a_1500_12478# 0.0187f
C213 w_n1594_38334# a_n1558_38434# 0.0187f
C214 a_1500_n3590# w_n1594_n3690# 0.0187f
C215 a_n1558_6298# a_n1558_5062# 0.0105f
C216 w_n1594_8670# a_n1500_9909# 0.0172f
C217 a_n1500_29685# a_n1500_28449# 3.11f
C218 w_n1594_4962# a_n1500_4965# 1.65f
C219 a_1500_n53030# w_n1594_n51894# 0.0023f
C220 a_n1558_n13478# a_n1558_n14714# 0.0105f
C221 a_n1500_n28407# a_1500_n28310# 0.217f
C222 w_n1594_18558# a_n1558_19894# 0.0023f
C223 a_n1558_58210# a_n1558_56974# 0.0105f
C224 a_n1558_13714# a_n1558_14950# 0.0105f
C225 a_1500_14950# a_1500_16186# 0.0105f
C226 a_n1500_50697# a_n1500_49461# 3.11f
C227 w_n1594_46986# a_n1500_48225# 0.0172f
C228 a_1500_n9770# a_n1500_n9867# 0.217f
C229 a_n1500_18561# a_n1500_17325# 3.11f
C230 a_n1500_n37059# a_n1500_n38295# 3.11f
C231 a_1500_n17186# a_1500_n15950# 0.0105f
C232 a_1500_n24602# w_n1594_n23466# 0.0023f
C233 a_n1558_27310# a_n1558_28546# 0.0105f
C234 a_n1500_29685# w_n1594_30918# 0.0172f
C235 w_n1594_n39534# a_1500_n40670# 0.0023f
C236 a_n1558_34726# w_n1594_34626# 0.0187f
C237 a_n1500_45753# a_1500_45850# 0.217f
C238 a_n1558_n56738# a_n1558_n57974# 0.0105f
C239 a_n1558_n8534# a_n1558_n9770# 0.0105f
C240 a_n1558_60682# a_n1558_59446# 0.0105f
C241 a_n1500_23505# a_1500_23602# 0.217f
C242 a_1500_n1118# a_1500_118# 0.0105f
C243 w_n1594_49458# a_n1500_49461# 1.65f
C244 a_n1500_n55599# a_1500_n55502# 0.217f
C245 w_n1594_n42006# a_n1558_n41906# 0.0187f
C246 a_n1558_53266# w_n1594_51930# 0.0023f
C247 w_n1594_n13578# a_n1558_n14714# 0.0023f
C248 w_n1594_2490# a_n1558_2590# 0.0187f
C249 a_1500_53266# w_n1594_53166# 0.0187f
C250 a_n1558_n53030# a_n1558_n54266# 0.0105f
C251 a_n1500_28449# a_n1558_28546# 0.217f
C252 a_n1558_23602# w_n1594_23502# 0.0187f
C253 w_n1594_n28410# a_n1500_n28407# 1.65f
C254 a_n1558_26074# w_n1594_27210# 0.0023f
C255 a_n1500_2493# a_1500_2590# 0.217f
C256 a_n1500_27213# a_1500_27310# 0.217f
C257 a_n1500_21# a_n1500_n1215# 3.11f
C258 a_1500_28546# a_n1500_28449# 0.217f
C259 a_n1558_n48086# w_n1594_n49422# 0.0023f
C260 a_1500_21130# w_n1594_22266# 0.0023f
C261 a_n1558_n53030# w_n1594_n53130# 0.0187f
C262 a_n1500_n38295# a_n1500_n39531# 3.11f
C263 w_n1594_13614# a_n1500_14853# 0.0172f
C264 w_n1594_4962# a_1500_5062# 0.0187f
C265 a_n1500_56877# w_n1594_58110# 0.0172f
C266 w_n1594_7434# a_n1500_8673# 0.0172f
C267 a_n1500_n12339# a_n1558_n12242# 0.217f
C268 w_n1594_17322# a_1500_18658# 0.0023f
C269 a_n1500_50697# a_n1500_51933# 3.11f
C270 w_n1594_n63018# a_n1500_n63015# 1.65f
C271 a_n1500_33393# a_1500_33490# 0.217f
C272 a_n1558_16186# a_n1558_14950# 0.0105f
C273 a_n1558_n53030# w_n1594_n54366# 0.0023f
C274 a_n1558_n2354# a_n1558_n1118# 0.0105f
C275 a_1500_n46850# w_n1594_n46950# 0.0187f
C276 a_n1558_3826# w_n1594_2490# 0.0023f
C277 a_1500_31018# a_1500_32254# 0.0105f
C278 a_1500_14950# w_n1594_16086# 0.0023f
C279 a_n1500_n24699# a_n1500_n23463# 3.11f
C280 a_n1558_53266# w_n1594_54402# 0.0023f
C281 a_n1500_n42003# a_1500_n41906# 0.217f
C282 a_n1558_n4826# a_n1558_n3590# 0.0105f
C283 w_n1594_n37062# a_1500_n36962# 0.0187f
C284 w_n1594_n18522# a_n1558_n18422# 0.0187f
C285 a_n1558_13714# w_n1594_13614# 0.0187f
C286 w_n1594_n35826# a_1500_n34490# 0.0023f
C287 a_n1500_1257# w_n1594_2490# 0.0172f
C288 a_n1558_50794# w_n1594_51930# 0.0023f
C289 a_n1500_56877# a_1500_56974# 0.217f
C290 w_n1594_n1218# a_n1558_n1118# 0.0187f
C291 w_n1594_n58074# a_1500_n59210# 0.0023f
C292 a_1500_n2354# w_n1594_n3690# 0.0023f
C293 a_1500_n48086# w_n1594_n48186# 0.0187f
C294 w_n1594_n27174# a_n1558_n27074# 0.0187f
C295 a_1500_37198# w_n1594_37098# 0.0187f
C296 a_n1500_n18519# a_n1500_n17283# 3.11f
C297 a_1500_n51794# w_n1594_n51894# 0.0187f
C298 a_1500_n23366# w_n1594_n22230# 0.0023f
C299 a_1500_59446# a_n1500_59349# 0.217f
C300 w_n1594_n35826# a_1500_n36962# 0.0023f
C301 a_n1558_n27074# a_n1558_n28310# 0.0105f
C302 w_n1594_46986# a_1500_47086# 0.0187f
C303 w_n1594_n2454# a_n1500_n1215# 0.0172f
C304 a_n1558_42142# w_n1594_42042# 0.0187f
C305 a_n1500_n23463# a_n1500_n22227# 3.11f
C306 w_n1594_n59310# a_1500_n60446# 0.0023f
C307 w_n1594_30918# a_n1558_31018# 0.0187f
C308 a_n1500_n49419# a_n1500_n50655# 3.11f
C309 a_1500_n51794# w_n1594_n50658# 0.0023f
C310 w_n1594_24738# a_1500_23602# 0.0023f
C311 a_1500_n23366# w_n1594_n23466# 0.0187f
C312 w_n1594_12378# a_n1500_11145# 0.0172f
C313 a_n1500_14853# w_n1594_14850# 1.65f
C314 w_n1594_n39534# a_1500_n39434# 0.0187f
C315 a_n1500_n14811# w_n1594_n13578# 0.0172f
C316 a_n1500_59349# a_n1558_59446# 0.217f
C317 a_n1500_n56835# a_1500_n56738# 0.217f
C318 a_n1500_n25935# a_n1500_n27171# 3.11f
C319 a_n1558_38434# a_n1500_38337# 0.217f
C320 w_n1594_45750# a_n1558_44614# 0.0023f
C321 a_n1558_27310# a_n1558_26074# 0.0105f
C322 a_n1558_61918# a_n1558_60682# 0.0105f
C323 w_n1594_n42006# a_n1558_n40670# 0.0023f
C324 a_n1500_n17283# w_n1594_n17286# 1.65f
C325 a_n1500_n53127# a_1500_n53030# 0.217f
C326 a_1500_37198# w_n1594_35862# 0.0023f
C327 w_n1594_n19758# a_n1500_n19755# 1.65f
C328 w_n1594_n12342# a_1500_n12242# 0.0187f
C329 w_n1594_9906# a_n1558_10006# 0.0187f
C330 a_n1558_13714# w_n1594_14850# 0.0023f
C331 w_n1594_29682# a_n1500_30921# 0.0172f
C332 a_1500_n59210# a_1500_n60446# 0.0105f
C333 a_n1500_n60543# a_n1558_n60446# 0.217f
C334 a_n1558_n51794# w_n1594_n53130# 0.0023f
C335 w_n1594_45750# a_n1500_46989# 0.0172f
C336 a_n1558_54502# a_n1500_54405# 0.217f
C337 a_n1500_7437# a_1500_7534# 0.217f
C338 w_n1594_32154# a_n1558_31018# 0.0023f
C339 a_n1558_n9770# w_n1594_n9870# 0.0187f
C340 w_n1594_n63018# a_n1500_n61779# 0.0172f
C341 a_1500_n30782# w_n1594_n29646# 0.0023f
C342 a_n1558_n23366# a_n1558_n22130# 0.0105f
C343 w_n1594_1254# a_n1500_21# 0.0172f
C344 w_n1594_3726# a_n1558_5062# 0.0023f
C345 a_1500_n45614# w_n1594_n46950# 0.0023f
C346 a_1500_24838# a_1500_26074# 0.0105f
C347 a_1500_39670# w_n1594_39570# 0.0187f
C348 w_n1594_28446# a_n1558_27310# 0.0023f
C349 a_n1500_n20991# a_n1500_n22227# 3.11f
C350 a_1500_21130# w_n1594_21030# 0.0187f
C351 a_n1558_n40670# a_n1558_n41906# 0.0105f
C352 a_1500_35962# a_1500_34726# 0.0105f
C353 a_n1500_n29643# a_n1500_n30879# 3.11f
C354 a_1500_26074# w_n1594_25974# 0.0187f
C355 a_1500_50794# a_1500_49558# 0.0105f
C356 w_n1594_19794# a_1500_18658# 0.0023f
C357 a_1500_53266# a_1500_54502# 0.0105f
C358 a_1500_n15950# a_n1500_n16047# 0.217f
C359 a_n1500_n32115# a_n1500_n33351# 3.11f
C360 w_n1594_28446# a_n1500_28449# 1.65f
C361 w_n1594_n58074# a_1500_n57974# 0.0187f
C362 a_1500_43378# w_n1594_42042# 0.0023f
C363 a_n1500_n34587# a_n1500_n35823# 3.11f
C364 a_n1500_n45711# a_n1558_n45614# 0.217f
C365 a_1500_n46850# w_n1594_n48186# 0.0023f
C366 a_1500_n44378# a_1500_n45614# 0.0105f
C367 a_n1500_22269# w_n1594_22266# 1.65f
C368 a_n1500_45753# w_n1594_44514# 0.0172f
C369 a_1500_n32018# w_n1594_n32118# 0.0187f
C370 a_1500_6298# w_n1594_7434# 0.0023f
C371 w_n1594_n22230# a_n1558_n22130# 0.0187f
C372 a_n1558_n20894# a_n1558_n22130# 0.0105f
C373 a_n1558_16186# w_n1594_14850# 0.0023f
C374 a_1500_38434# a_1500_39670# 0.0105f
C375 a_1500_n32018# w_n1594_n30882# 0.0023f
C376 a_n1500_6201# w_n1594_7434# 0.0172f
C377 a_n1500_43281# w_n1594_42042# 0.0172f
C378 a_n1500_55641# a_n1500_54405# 3.11f
C379 a_1500_n50558# w_n1594_n51894# 0.0023f
C380 a_n1500_n11103# w_n1594_n11106# 1.65f
C381 w_n1594_n19758# a_1500_n19658# 0.0187f
C382 w_n1594_37098# a_1500_35962# 0.0023f
C383 a_n1558_55738# w_n1594_56874# 0.0023f
C384 w_n1594_n40770# a_n1500_n42003# 0.0172f
C385 w_n1594_33390# a_n1558_33490# 0.0187f
C386 w_n1594_n59310# a_1500_n59210# 0.0187f
C387 a_n1558_10006# w_n1594_8670# 0.0023f
C388 a_n1558_n22130# w_n1594_n23466# 0.0023f
C389 a_1500_n50558# w_n1594_n50658# 0.0187f
C390 a_1500_3826# a_n1500_3729# 0.217f
C391 a_n1500_n23463# w_n1594_n24702# 0.0172f
C392 w_n1594_n39534# a_1500_n38198# 0.0023f
C393 a_n1558_32254# w_n1594_30918# 0.0023f
C394 a_1500_1354# w_n1594_1254# 0.0187f
C395 a_n1558_1354# w_n1594_18# 0.0023f
C396 a_n1558_16186# a_n1558_17422# 0.0105f
C397 a_n1558_n2354# a_n1558_n3590# 0.0105f
C398 a_n1500_n7395# w_n1594_n8634# 0.0172f
C399 a_n1558_34726# a_n1558_33490# 0.0105f
C400 a_1500_13714# w_n1594_12378# 0.0023f
C401 a_n1500_n17283# w_n1594_n16050# 0.0172f
C402 a_1500_n13478# w_n1594_n14814# 0.0023f
C403 a_1500_42142# w_n1594_42042# 0.0187f
C404 a_1500_n7298# a_1500_n8534# 0.0105f
C405 a_n1558_32254# a_n1500_32157# 0.217f
C406 a_n1558_n51794# a_n1558_n53030# 0.0105f
C407 a_n1500_n20991# a_n1500_n19755# 3.11f
C408 a_n1500_21033# a_n1500_19797# 3.11f
C409 a_1500_35962# w_n1594_35862# 0.0187f
C410 w_n1594_49458# a_n1558_48322# 0.0023f
C411 w_n1594_33390# a_n1500_33393# 1.65f
C412 a_n1558_n15950# w_n1594_n17286# 0.0023f
C413 w_n1594_39570# a_1500_40906# 0.0023f
C414 w_n1594_18558# a_1500_18658# 0.0187f
C415 a_1500_11242# a_1500_10006# 0.0105f
C416 w_n1594_n61782# a_n1558_n62918# 0.0023f
C417 a_n1500_21033# w_n1594_22266# 0.0172f
C418 a_1500_n29546# w_n1594_n29646# 0.0187f
C419 w_n1594_49458# a_1500_48322# 0.0023f
C420 a_n1500_n18519# w_n1594_n17286# 0.0172f
C421 a_n1500_n55599# w_n1594_n55602# 1.65f
C422 a_n1500_25977# a_1500_26074# 0.217f
C423 w_n1594_n13578# a_1500_n12242# 0.0023f
C424 a_n1558_32254# w_n1594_32154# 0.0187f
C425 a_1500_n20894# a_1500_n22130# 0.0105f
C426 a_n1500_n40767# a_1500_n40670# 0.217f
C427 a_1500_n45614# w_n1594_n44478# 0.0023f
C428 a_n1500_45753# a_n1500_46989# 3.11f
C429 w_n1594_50694# a_1500_49558# 0.0023f
C430 w_n1594_n58074# a_1500_n56738# 0.0023f
C431 a_n1500_n20991# w_n1594_n20994# 1.65f
C432 w_n1594_4962# a_n1500_3729# 0.0172f
C433 a_n1500_16089# w_n1594_14850# 0.0172f
C434 a_n1558_n32018# w_n1594_n33354# 0.0023f
C435 a_1500_118# a_n1500_21# 0.217f
C436 a_n1558_12478# w_n1594_12378# 0.0187f
C437 a_1500_n30782# w_n1594_n32118# 0.0023f
C438 w_n1594_3726# a_n1500_4965# 0.0172f
C439 w_n1594_n12342# a_n1558_n11006# 0.0023f
C440 w_n1594_n20994# a_1500_n20894# 0.0187f
C441 a_1500_n30782# w_n1594_n30882# 0.0187f
C442 a_n1558_40906# w_n1594_40806# 0.0187f
C443 a_n1558_n23366# w_n1594_n22230# 0.0023f
C444 a_1500_n8534# w_n1594_n7398# 0.0023f
C445 a_1500_8770# a_1500_10006# 0.0105f
C446 a_1500_54502# w_n1594_53166# 0.0023f
C447 a_1500_23602# a_1500_24838# 0.0105f
C448 w_n1594_n40770# a_n1500_n40767# 1.65f
C449 a_1500_n19658# a_1500_n20894# 0.0105f
C450 a_n1558_8770# a_n1500_8673# 0.217f
C451 a_1500_8770# a_1500_7534# 0.0105f
C452 a_1500_38434# w_n1594_37098# 0.0023f
C453 w_n1594_n59310# a_1500_n57974# 0.0023f
C454 a_n1500_n48183# a_n1500_n49419# 3.11f
C455 w_n1594_n28410# a_n1500_n27171# 0.0172f
C456 a_n1500_n24699# a_n1500_n25935# 3.11f
C457 a_n1558_n23366# w_n1594_n23466# 0.0187f
C458 a_n1500_21033# a_n1558_21130# 0.217f
C459 a_1500_6298# w_n1594_6198# 0.0187f
C460 w_n1594_16086# a_1500_16186# 0.0187f
C461 a_1500_n49322# w_n1594_n50658# 0.0023f
C462 a_n1500_22269# w_n1594_21030# 0.0172f
C463 w_n1594_13614# a_n1500_13617# 1.65f
C464 w_n1594_50694# a_n1558_49558# 0.0023f
C465 a_n1500_6201# w_n1594_6198# 1.65f
C466 a_n1500_n13575# a_1500_n13478# 0.217f
C467 a_n1500_1257# w_n1594_18# 0.0172f
C468 a_n1500_58113# w_n1594_56874# 0.0172f
C469 w_n1594_n22230# a_n1558_n20894# 0.0023f
C470 a_n1500_n51891# a_1500_n51794# 0.217f
C471 a_1500_34726# w_n1594_34626# 0.0187f
C472 a_n1558_45850# w_n1594_44514# 0.0023f
C473 a_n1558_n2354# w_n1594_n1218# 0.0023f
C474 a_n1558_48322# a_n1558_47086# 0.0105f
C475 a_1500_n44378# a_1500_n43142# 0.0105f
C476 w_n1594_60582# a_1500_60682# 0.0187f
C477 a_n1558_n44378# a_n1500_n44475# 0.217f
C478 w_n1594_11142# a_1500_10006# 0.0023f
C479 a_n1500_28449# w_n1594_29682# 0.0172f
C480 w_n1594_3726# a_1500_5062# 0.0023f
C481 a_1500_n57974# a_1500_n59210# 0.0105f
C482 a_n1558_n6062# w_n1594_n4926# 0.0023f
C483 a_n1500_n59307# a_n1558_n59210# 0.217f
C484 a_n1500_n8631# a_1500_n8534# 0.217f
C485 a_n1558_58210# w_n1594_59346# 0.0023f
C486 a_n1558_n15950# w_n1594_n14814# 0.0023f
C487 a_n1558_n19658# a_n1558_n20894# 0.0105f
C488 a_1500_n7298# w_n1594_n8634# 0.0023f
C489 w_n1594_n6162# a_n1558_n7298# 0.0023f
C490 a_n1558_61918# a_n1500_61821# 0.217f
C491 a_1500_1354# a_1500_118# 0.0105f
C492 a_n1558_n9770# a_n1558_n11006# 0.0105f
C493 a_n1558_n15950# w_n1594_n16050# 0.0187f
C494 a_n1558_23602# a_n1558_24838# 0.0105f
C495 w_n1594_n43242# a_n1500_n44475# 0.0172f
C496 w_n1594_45750# a_n1500_45753# 1.65f
C497 w_n1594_n61782# a_n1558_n61682# 0.0187f
C498 a_n1500_n55599# a_n1558_n55502# 0.217f
C499 a_n1558_53266# a_n1558_52030# 0.0105f
C500 a_n1558_43378# w_n1594_42042# 0.0023f
C501 w_n1594_n27174# a_n1558_n25838# 0.0023f
C502 w_n1594_n25938# a_n1500_n27171# 0.0172f
C503 a_n1558_3826# a_n1500_3729# 0.217f
C504 a_n1558_118# a_n1500_21# 0.217f
C505 a_n1558_53266# a_n1500_53169# 0.217f
C506 a_n1500_n46947# w_n1594_n45714# 0.0172f
C507 a_n1500_n54363# w_n1594_n55602# 0.0172f
C508 w_n1594_11142# a_n1558_11242# 0.0187f
C509 a_n1558_n39434# a_n1558_n40670# 0.0105f
C510 a_1500_n44378# w_n1594_n44478# 0.0187f
C511 a_n1500_18561# a_n1500_19797# 3.11f
C512 a_1500_n27074# a_n1500_n27171# 0.217f
C513 a_n1500_21033# w_n1594_21030# 1.65f
C514 a_n1500_13617# w_n1594_14850# 0.0172f
C515 w_n1594_n60546# a_n1558_n61682# 0.0023f
C516 a_1500_43378# w_n1594_44514# 0.0023f
C517 a_n1500_n33351# a_n1500_n34587# 3.11f
C518 w_n1594_n38298# a_n1500_n37059# 0.0172f
C519 a_n1500_23505# a_n1500_24741# 3.11f
C520 a_n1500_n55599# w_n1594_n56838# 0.0172f
C521 w_n1594_n34590# a_n1558_n35726# 0.0023f
C522 a_n1558_45850# a_n1558_44614# 0.0105f
C523 a_n1500_39573# a_1500_39670# 0.217f
C524 a_n1500_42045# w_n1594_40806# 0.0172f
C525 a_1500_n29546# w_n1594_n30882# 0.0023f
C526 a_n1500_43281# w_n1594_44514# 0.0172f
C527 a_n1500_n32115# a_1500_n32018# 0.217f
C528 a_n1500_29685# a_1500_29782# 0.217f
C529 a_n1558_n29546# a_n1558_n28310# 0.0105f
C530 a_n1558_n8534# w_n1594_n8634# 0.0187f
C531 w_n1594_n40770# a_n1500_n39531# 0.0172f
C532 a_n1558_52030# a_n1558_50794# 0.0105f
C533 a_n1500_n6159# a_n1558_n6062# 0.217f
C534 a_n1500_37101# w_n1594_37098# 1.65f
C535 a_1500_n6062# w_n1594_n6162# 0.0187f
C536 a_1500_40906# a_n1500_40809# 0.217f
C537 a_1500_27310# w_n1594_25974# 0.0023f
C538 w_n1594_48222# a_n1558_47086# 0.0023f
C539 w_n1594_24738# a_n1500_23505# 0.0172f
C540 a_1500_39670# w_n1594_38334# 0.0023f
C541 a_n1500_12381# w_n1594_13614# 0.0172f
C542 a_1500_21130# w_n1594_19794# 0.0023f
C543 a_1500_n13478# a_1500_n14714# 0.0105f
C544 a_n1500_n18519# a_n1500_n19755# 3.11f
C545 w_n1594_n38298# a_n1500_n39531# 0.0172f
C546 a_1500_n8534# w_n1594_n9870# 0.0023f
C547 a_n1500_11145# a_n1558_11242# 0.217f
C548 a_n1500_48225# a_n1500_49461# 3.11f
C549 a_n1558_12478# a_n1558_13714# 0.0105f
C550 a_n1558_n9770# a_n1500_n9867# 0.217f
C551 w_n1594_n44478# a_1500_n43142# 0.0023f
C552 a_n1500_n4923# a_n1500_n3687# 3.11f
C553 a_n1558_n50558# a_n1558_n51794# 0.0105f
C554 a_1500_14950# a_n1500_14853# 0.217f
C555 a_n1500_n29643# w_n1594_n28410# 0.0172f
C556 a_n1558_n4826# w_n1594_n4926# 0.0187f
C557 a_1500_44614# a_1500_45850# 0.0105f
C558 a_1500_23602# w_n1594_23502# 0.0187f
C559 w_n1594_n18522# a_n1500_n17283# 0.0172f
C560 w_n1594_4962# a_1500_3826# 0.0023f
C561 a_n1500_37101# w_n1594_35862# 0.0172f
C562 w_n1594_16086# a_n1500_17325# 0.0172f
C563 a_1500_28546# a_1500_29782# 0.0105f
C564 a_n1558_40906# a_n1558_42142# 0.0105f
C565 a_1500_n9770# a_1500_n8534# 0.0105f
C566 w_n1594_56874# a_n1500_55641# 0.0172f
C567 w_n1594_n43242# a_n1500_n43239# 1.65f
C568 w_n1594_n61782# a_n1558_n60446# 0.0023f
C569 a_n1500_n1215# a_n1558_n1118# 0.217f
C570 a_1500_40906# w_n1594_42042# 0.0023f
C571 w_n1594_n55602# a_n1500_n56835# 0.0172f
C572 a_n1500_n8631# w_n1594_n8634# 1.65f
C573 w_n1594_n25938# a_n1500_n25935# 1.65f
C574 w_n1594_n37062# a_n1558_n36962# 0.0187f
C575 w_n1594_37098# a_n1500_35865# 0.0172f
C576 a_n1500_n25935# w_n1594_n24702# 0.0172f
C577 a_n1500_n45711# w_n1594_n45714# 1.65f
C578 a_n1500_12381# a_1500_12478# 0.217f
C579 a_n1500_n50655# w_n1594_n49422# 0.0172f
C580 w_n1594_59346# a_1500_59446# 0.0187f
C581 a_1500_58210# w_n1594_59346# 0.0023f
C582 a_n1500_n61779# a_n1500_n63015# 3.11f
C583 a_n1500_n39531# a_1500_n39434# 0.217f
C584 w_n1594_24738# a_n1500_24741# 1.65f
C585 w_n1594_49458# a_1500_49558# 0.0187f
C586 w_n1594_54402# a_1500_55738# 0.0023f
C587 a_n1558_n27074# a_n1558_n25838# 0.0105f
C588 a_1500_n11006# w_n1594_n9870# 0.0023f
C589 a_n1558_34726# a_n1558_35962# 0.0105f
C590 w_n1594_17322# a_n1558_17422# 0.0187f
C591 a_n1500_n4923# w_n1594_n6162# 0.0172f
C592 w_n1594_n56838# a_n1500_n58071# 0.0172f
C593 a_n1558_54502# w_n1594_53166# 0.0023f
C594 a_n1558_18658# a_n1558_19894# 0.0105f
C595 a_n1500_n55599# w_n1594_n54366# 0.0172f
C596 w_n1594_n60546# a_n1558_n60446# 0.0187f
C597 w_n1594_n29646# a_n1558_n28310# 0.0023f
C598 w_n1594_46986# a_n1558_48322# 0.0023f
C599 a_n1500_37101# a_n1558_37198# 0.217f
C600 w_n1594_n34590# a_n1558_n34490# 0.0187f
C601 w_n1594_59346# a_n1558_59446# 0.0187f
C602 w_n1594_n33354# a_n1558_n34490# 0.0023f
C603 a_n1500_29685# a_n1558_29782# 0.217f
C604 a_n1500_n43239# a_n1558_n43142# 0.217f
C605 w_n1594_n4926# a_n1558_n3590# 0.0023f
C606 w_n1594_55638# a_1500_55738# 0.0187f
C607 a_1500_n41906# a_1500_n43142# 0.0105f
C608 a_n1500_7437# a_n1558_7534# 0.217f
C609 a_n1500_n2451# a_n1500_n3687# 3.11f
C610 w_n1594_n32118# a_1500_n33254# 0.0023f
C611 w_n1594_n35826# a_n1558_n36962# 0.0023f
C612 w_n1594_45750# a_n1558_45850# 0.0187f
C613 w_n1594_56874# a_n1558_56974# 0.0187f
C614 a_n1558_n30782# a_n1558_n32018# 0.0105f
C615 a_n1500_35865# w_n1594_35862# 1.65f
C616 a_n1558_n4826# w_n1594_n3690# 0.0023f
C617 a_n1558_n35726# a_n1558_n36962# 0.0105f
C618 a_1500_n11006# a_1500_n9770# 0.0105f
C619 a_n1500_n46947# a_n1500_n48183# 3.11f
C620 w_n1594_46986# a_1500_48322# 0.0023f
C621 a_n1500_n11103# a_n1500_n12339# 3.11f
C622 w_n1594_n45714# a_n1500_n44475# 0.0172f
C623 w_n1594_49458# a_n1558_49558# 0.0187f
C624 w_n1594_n38298# a_n1500_n38295# 1.65f
C625 w_n1594_n11106# a_n1500_n12339# 0.0172f
C626 a_1500_28546# a_1500_27310# 0.0105f
C627 a_1500_n11006# a_1500_n12242# 0.0105f
C628 a_n1500_27213# w_n1594_25974# 0.0172f
C629 a_n1558_28546# a_n1558_29782# 0.0105f
C630 a_1500_10006# a_n1500_9909# 0.217f
C631 a_n1558_n6062# w_n1594_n7398# 0.0023f
C632 a_n1500_n50655# a_1500_n50558# 0.217f
C633 w_n1594_18# a_n1500_n1215# 0.0172f
C634 a_n1500_51933# w_n1594_51930# 1.65f
C635 a_1500_31018# w_n1594_29682# 0.0023f
C636 a_n1500_34629# w_n1594_34626# 1.65f
C637 w_n1594_17322# a_1500_17422# 0.0187f
C638 w_n1594_2490# a_n1500_2493# 1.65f
C639 a_n1558_n36962# a_n1558_n38198# 0.0105f
C640 a_n1500_12381# w_n1594_11142# 0.0172f
C641 a_1500_n1118# w_n1594_n2454# 0.0023f
C642 a_n1558_8770# a_n1558_10006# 0.0105f
C643 a_1500_1354# a_1500_2590# 0.0105f
C644 a_n1558_1354# a_n1558_2590# 0.0105f
C645 a_n1500_n24699# w_n1594_n25938# 0.0172f
C646 a_n1500_n58071# a_n1558_n57974# 0.217f
C647 a_1500_n56738# a_1500_n57974# 0.0105f
C648 a_n1558_32254# a_n1558_33490# 0.0105f
C649 a_n1500_42045# a_n1558_42142# 0.217f
C650 a_n1500_n24699# w_n1594_n24702# 1.65f
C651 a_n1500_44517# w_n1594_44514# 1.65f
C652 w_n1594_n43242# a_n1500_n42003# 0.0172f
C653 w_n1594_n42006# a_n1500_n43239# 0.0172f
C654 a_1500_n53030# a_1500_n54266# 0.0105f
C655 a_n1500_n54363# a_n1558_n54266# 0.217f
C656 a_n1558_42142# w_n1594_40806# 0.0023f
C657 w_n1594_30918# a_n1500_30921# 1.65f
C658 a_n1500_6201# a_n1500_4965# 3.11f
C659 a_n1558_43378# w_n1594_44514# 0.0023f
C660 w_n1594_n28410# a_1500_n28310# 0.0187f
C661 w_n1594_n37062# a_n1558_n35726# 0.0023f
C662 w_n1594_33390# a_1500_33490# 0.0187f
C663 a_n1558_n3590# w_n1594_n3690# 0.0187f
C664 a_1500_n9770# w_n1594_n8634# 0.0023f
C665 a_n1500_n49419# w_n1594_n49422# 1.65f
C666 a_n1500_32157# a_n1500_30921# 3.11f
C667 w_n1594_60582# a_n1558_60682# 0.0187f
C668 a_n1500_n22227# a_1500_n22130# 0.217f
C669 a_n1500_n54363# w_n1594_n53130# 0.0172f
C670 w_n1594_n18522# a_n1500_n18519# 1.65f
C671 a_n1558_n38198# a_n1558_n39434# 0.0105f
C672 w_n1594_61818# a_n1558_61918# 0.0187f
C673 a_n1558_n11006# a_n1558_n12242# 0.0105f
C674 a_n1558_6298# a_n1558_7534# 0.0105f
C675 a_n1500_56877# w_n1594_56874# 1.65f
C676 a_1500_32254# a_1500_33490# 0.0105f
C677 a_n1558_29782# a_n1558_31018# 0.0105f
C678 a_n1500_n13575# w_n1594_n14814# 0.0172f
C679 w_n1594_n63018# a_1500_n62918# 0.0187f
C680 w_n1594_n12342# a_n1558_n13478# 0.0023f
C681 a_n1558_23602# a_n1558_22366# 0.0105f
C682 a_1500_n2354# a_1500_n1118# 0.0105f
C683 w_n1594_3726# a_n1500_3729# 1.65f
C684 w_n1594_55638# a_1500_56974# 0.0023f
C685 w_n1594_n56838# a_n1500_n56835# 1.65f
C686 a_n1558_44614# w_n1594_43278# 0.0023f
C687 w_n1594_28446# a_1500_29782# 0.0023f
C688 a_n1500_n54363# w_n1594_n54366# 1.65f
C689 w_n1594_n60546# a_n1558_n59210# 0.0023f
C690 a_1500_17422# a_1500_18658# 0.0105f
C691 a_n1558_n48086# w_n1594_n46950# 0.0023f
C692 a_n1500_1257# a_n1558_1354# 0.217f
C693 a_n1558_3826# w_n1594_4962# 0.0023f
C694 w_n1594_n34590# a_n1558_n33254# 0.0023f
C695 w_n1594_n20994# a_n1500_n22227# 0.0172f
C696 a_n1558_n24602# a_n1558_n23366# 0.0105f
C697 w_n1594_n33354# a_n1558_n33254# 0.0187f
C698 a_1500_37198# a_1500_35962# 0.0105f
C699 w_n1594_n37062# a_n1558_n38198# 0.0023f
C700 a_n1558_12478# a_n1558_11242# 0.0105f
C701 a_n1500_12381# a_n1500_11145# 3.11f
C702 w_n1594_n35826# a_n1558_n35726# 0.0187f
C703 a_n1500_n30879# a_1500_n30782# 0.217f
C704 w_n1594_46986# a_1500_45850# 0.0023f
C705 a_n1500_22269# a_n1500_23505# 3.11f
C706 a_n1558_52030# w_n1594_51930# 0.0187f
C707 a_1500_6298# a_1500_5062# 0.0105f
C708 w_n1594_32154# a_n1500_30921# 0.0172f
C709 a_1500_44614# w_n1594_44514# 0.0187f
C710 a_1500_13714# a_n1500_13617# 0.217f
C711 a_n1500_53169# w_n1594_51930# 0.0172f
C712 a_n1558_37198# w_n1594_38334# 0.0023f
C713 a_n1500_n35823# a_1500_n35726# 0.217f
C714 w_n1594_n27174# a_n1500_n28407# 0.0172f
C715 a_n1558_n49322# w_n1594_n48186# 0.0023f
C716 a_n1500_44517# a_n1558_44614# 0.217f
C717 a_n1558_55738# a_n1558_54502# 0.0105f
C718 a_n1558_27310# w_n1594_27210# 0.0187f
C719 a_n1500_27213# a_n1500_25977# 3.11f
C720 a_n1558_43378# a_n1558_44614# 0.0105f
C721 w_n1594_n4926# a_1500_n4826# 0.0187f
C722 a_n1558_45850# a_n1500_45753# 0.217f
C723 a_n1558_n53030# w_n1594_n51894# 0.0023f
C724 a_1500_52030# w_n1594_51930# 0.0187f
C725 a_1500_n27074# a_1500_n28310# 0.0105f
C726 a_n1500_28449# w_n1594_27210# 0.0172f
C727 a_1500_n3590# a_n1500_n3687# 0.217f
C728 a_n1500_n28407# a_n1558_n28310# 0.217f
C729 w_n1594_50694# a_1500_50794# 0.0187f
C730 a_n1500_21033# w_n1594_19794# 0.0172f
C731 a_n1500_34629# a_n1500_35865# 3.11f
C732 a_n1558_n49322# a_n1558_n50558# 0.0105f
C733 a_n1558_3826# a_n1558_2590# 0.0105f
C734 a_n1500_48225# a_n1558_48322# 0.217f
C735 a_n1558_8770# w_n1594_9906# 0.0023f
C736 a_n1500_43281# a_n1500_42045# 3.11f
C737 a_n1500_n37059# a_1500_n36962# 0.217f
C738 w_n1594_4962# a_n1558_6298# 0.0023f
C739 a_n1558_n24602# w_n1594_n23466# 0.0023f
C740 w_n1594_17322# a_n1500_18561# 0.0172f
C741 w_n1594_n39534# a_n1558_n40670# 0.0023f
C742 w_n1594_n19758# a_1500_n18422# 0.0023f
C743 w_n1594_54402# a_n1500_53169# 0.0172f
C744 a_1500_n54266# a_1500_n55502# 0.0105f
C745 a_n1558_n15950# a_n1558_n14714# 0.0105f
C746 w_n1594_n42006# a_n1500_n42003# 1.65f
C747 a_n1558_n2354# w_n1594_n3690# 0.0023f
C748 a_n1558_55738# a_n1500_55641# 0.217f
C749 a_1500_48322# a_n1500_48225# 0.217f
C750 w_n1594_n20994# a_n1500_n19755# 0.0172f
C751 w_n1594_n28410# a_1500_n27074# 0.0023f
C752 a_n1500_24741# a_1500_24838# 0.217f
C753 a_1500_6298# a_1500_7534# 0.0105f
C754 w_n1594_28446# a_1500_27310# 0.0023f
C755 a_n1500_n48183# w_n1594_n49422# 0.0172f
C756 w_n1594_60582# a_n1500_59349# 0.0172f
C757 w_n1594_37098# a_n1500_38337# 0.0172f
C758 a_n1500_n17283# a_1500_n17186# 0.217f
C759 a_n1500_n60543# a_n1500_n61779# 3.11f
C760 a_n1500_n53127# w_n1594_n53130# 1.65f
C761 a_n1500_n38295# a_1500_n38198# 0.217f
C762 a_n1500_42045# a_1500_42142# 0.217f
C763 a_1500_n19658# a_n1500_n19755# 0.217f
C764 a_1500_n14714# w_n1594_n14814# 0.0187f
C765 a_n1500_24741# w_n1594_25974# 0.0172f
C766 w_n1594_28446# a_n1558_29782# 0.0023f
C767 a_n1500_n2451# w_n1594_n2454# 1.65f
C768 w_n1594_n63018# a_1500_n61682# 0.0023f
C769 w_n1594_n16050# a_1500_n14714# 0.0023f
C770 a_1500_42142# w_n1594_40806# 0.0023f
C771 w_n1594_18558# a_n1558_17422# 0.0023f
C772 a_n1558_n19658# a_n1558_n18422# 0.0105f
C773 w_n1594_17322# a_n1558_18658# 0.0023f
C774 a_n1500_n53127# w_n1594_n54366# 0.0172f
C775 a_1500_n4826# w_n1594_n3690# 0.0023f
C776 w_n1594_24738# a_1500_24838# 0.0187f
C777 a_n1500_n3687# w_n1594_n2454# 0.0172f
C778 w_n1594_n20994# a_1500_n22130# 0.0023f
C779 a_n1558_n46850# w_n1594_n46950# 0.0187f
C780 a_1500_56974# a_1500_55738# 0.0105f
C781 a_n1558_n18422# a_n1558_n17186# 0.0105f
C782 a_1500_n23366# a_n1500_n23463# 0.217f
C783 w_n1594_13614# a_n1558_14950# 0.0023f
C784 a_n1500_18561# a_1500_18658# 0.217f
C785 a_n1500_n42003# a_n1558_n41906# 0.217f
C786 a_1500_n40670# a_1500_n41906# 0.0105f
C787 w_n1594_n35826# a_n1558_n34490# 0.0023f
C788 a_n1558_n29546# a_n1558_n30782# 0.0105f
C789 a_1500_38434# a_1500_37198# 0.0105f
C790 a_n1500_46989# a_n1558_47086# 0.217f
C791 a_n1558_55738# a_n1558_56974# 0.0105f
C792 a_n1558_n32018# a_n1558_n33254# 0.0105f
C793 w_n1594_n13578# a_n1558_n13478# 0.0187f
C794 a_n1558_8770# w_n1594_8670# 0.0187f
C795 w_n1594_48222# a_n1500_48225# 1.65f
C796 w_n1594_n58074# a_n1558_n59210# 0.0023f
C797 a_n1558_n34490# a_n1558_n35726# 0.0105f
C798 a_n1558_n48086# w_n1594_n48186# 0.0187f
C799 w_n1594_n25938# a_1500_n27074# 0.0023f
C800 a_n1500_n45711# a_n1500_n46947# 3.11f
C801 a_1500_n2354# a_n1500_n2451# 0.217f
C802 w_n1594_45750# a_n1500_44517# 0.0172f
C803 a_n1558_n51794# w_n1594_n51894# 0.0187f
C804 a_1500_n19658# w_n1594_n20994# 0.0023f
C805 a_n1558_n7298# w_n1594_n8634# 0.0023f
C806 a_1500_31018# a_n1500_30921# 0.217f
C807 w_n1594_2490# a_1500_2590# 0.0187f
C808 w_n1594_n40770# a_1500_n41906# 0.0023f
C809 w_n1594_n59310# a_n1558_n60446# 0.0023f
C810 a_n1500_n49419# a_1500_n49322# 0.217f
C811 a_1500_17422# w_n1594_18558# 0.0023f
C812 w_n1594_n1218# a_n1500_n1215# 1.65f
C813 a_n1500_23505# w_n1594_23502# 1.65f
C814 a_n1558_n51794# w_n1594_n50658# 0.0023f
C815 w_n1594_16086# a_n1500_14853# 0.0172f
C816 w_n1594_3726# a_1500_3826# 0.0187f
C817 w_n1594_n39534# a_n1558_n39434# 0.0187f
C818 a_1500_29782# w_n1594_29682# 0.0187f
C819 a_1500_n55502# a_1500_n56738# 0.0105f
C820 a_n1500_n56835# a_n1558_n56738# 0.217f
C821 a_n1500_n25935# a_1500_n25838# 0.217f
C822 a_n1558_58210# w_n1594_58110# 0.0187f
C823 w_n1594_58110# a_1500_56974# 0.0023f
C824 a_n1500_n12339# a_n1500_n13575# 3.11f
C825 w_n1594_n42006# a_n1500_n40767# 0.0172f
C826 a_1500_n51794# a_1500_n53030# 0.0105f
C827 a_n1500_n53127# a_n1558_n53030# 0.217f
C828 a_1500_48322# a_1500_47086# 0.0105f
C829 w_n1594_14850# a_n1558_14950# 0.0187f
C830 w_n1594_n18522# a_n1500_n19755# 0.0172f
C831 w_n1594_n12342# a_n1558_n12242# 0.0187f
C832 a_n1500_18561# w_n1594_19794# 0.0172f
C833 a_n1500_42045# w_n1594_43278# 0.0172f
C834 w_n1594_33390# a_1500_32254# 0.0023f
C835 a_n1500_25977# a_n1500_24741# 3.11f
C836 a_n1558_12478# a_n1500_12381# 0.217f
C837 a_1500_44614# w_n1594_45750# 0.0023f
C838 a_n1558_34726# w_n1594_33390# 0.0023f
C839 a_n1558_10006# a_n1558_11242# 0.0105f
C840 a_1500_n12242# a_1500_n13478# 0.0105f
C841 a_n1500_n51891# w_n1594_n53130# 0.0172f
C842 a_n1500_34629# a_n1500_33393# 3.11f
C843 w_n1594_28446# a_n1500_27213# 0.0172f
C844 a_n1558_49558# a_n1558_50794# 0.0105f
C845 a_n1558_n30782# w_n1594_n29646# 0.0023f
C846 a_n1558_118# a_n1558_n1118# 0.0105f
C847 w_n1594_45750# a_n1558_47086# 0.0023f
C848 a_n1558_8770# w_n1594_7434# 0.0023f
C849 w_n1594_18# a_1500_118# 0.0187f
C850 a_n1558_n45614# w_n1594_n46950# 0.0023f
C851 a_n1500_32157# w_n1594_30918# 0.0172f
C852 w_n1594_60582# a_n1500_61821# 0.0172f
C853 w_n1594_24738# a_n1500_25977# 0.0172f
C854 a_n1558_n14714# w_n1594_n14814# 0.0187f
C855 a_n1500_21033# a_1500_21130# 0.217f
C856 a_n1500_n29643# a_1500_n29546# 0.217f
C857 a_n1500_37101# a_1500_37198# 0.217f
C858 w_n1594_n16050# a_n1558_n14714# 0.0023f
C859 a_n1500_24741# w_n1594_23502# 0.0172f
C860 a_n1500_58113# a_n1500_59349# 3.11f
C861 w_n1594_48222# a_1500_47086# 0.0023f
C862 a_n1558_18658# w_n1594_19794# 0.0023f
C863 a_n1500_n9867# w_n1594_n8634# 0.0172f
C864 w_n1594_n58074# a_n1558_n57974# 0.0187f
C865 a_n1500_n34587# a_1500_n34490# 0.217f
C866 w_n1594_54402# a_n1500_54405# 1.65f
C867 a_1500_n3590# w_n1594_n2454# 0.0023f
C868 w_n1594_13614# a_1500_12478# 0.0023f
C869 a_n1558_n46850# w_n1594_n48186# 0.0023f
C870 a_n1500_50697# a_1500_50794# 0.217f
C871 a_n1558_n32018# w_n1594_n32118# 0.0187f
C872 a_n1558_n32018# w_n1594_n30882# 0.0023f
C873 w_n1594_16086# a_n1558_16186# 0.0187f
C874 a_n1558_n50558# w_n1594_n51894# 0.0023f
C875 w_n1594_55638# a_n1500_54405# 0.0172f
C876 a_1500_39670# w_n1594_40806# 0.0023f
C877 w_n1594_37098# a_n1558_35962# 0.0023f
C878 w_n1594_n18522# a_1500_n19658# 0.0023f
C879 w_n1594_n40770# a_1500_n40670# 0.0187f
C880 w_n1594_n59310# a_n1558_n59210# 0.0187f
C881 w_n1594_49458# a_1500_50794# 0.0023f
C882 a_n1558_n48086# a_n1558_n49322# 0.0105f
C883 a_n1500_n17283# a_n1500_n16047# 3.11f
C884 w_n1594_32154# a_n1500_32157# 1.65f
C885 a_n1558_n50558# w_n1594_n50658# 0.0187f
C886 a_n1558_n24602# a_n1558_n25838# 0.0105f
C887 a_1500_n17186# w_n1594_n17286# 0.0187f
C888 a_n1500_44517# a_n1500_45753# 3.11f
C889 w_n1594_29682# a_n1558_29782# 0.0187f
C890 a_n1500_n11103# w_n1594_n9870# 0.0172f
C891 a_n1500_2493# a_n1500_3729# 3.11f
C892 w_n1594_9906# a_1500_10006# 0.0187f
C893 a_n1500_18561# w_n1594_18558# 1.65f
C894 w_n1594_n39534# a_n1558_n38198# 0.0023f
C895 a_1500_11242# a_1500_12478# 0.0105f
C896 a_n1500_16089# a_1500_16186# 0.217f
C897 a_1500_47086# a_1500_45850# 0.0105f
C898 a_n1558_n6062# a_n1558_n7298# 0.0105f
C899 a_1500_61918# a_1500_60682# 0.0105f
C900 w_n1594_46986# a_n1500_46989# 1.65f
C901 a_1500_n2354# a_1500_n3590# 0.0105f
C902 w_n1594_3726# a_n1558_2590# 0.0023f
C903 a_n1558_53266# w_n1594_53166# 0.0187f
C904 w_n1594_18# a_n1558_118# 0.0187f
C905 a_n1500_51933# a_n1558_52030# 0.217f
C906 a_n1558_n12242# a_n1558_n13478# 0.0105f
C907 a_1500_35962# w_n1594_34626# 0.0023f
C908 a_n1558_35962# w_n1594_35862# 0.0187f
C909 a_n1500_51933# a_n1500_53169# 3.11f
C910 w_n1594_9906# a_n1558_11242# 0.0023f
C911 a_n1500_n45711# a_n1500_n44475# 3.11f
C912 a_n1558_22366# w_n1594_22266# 0.0187f
C913 a_1500_n11006# w_n1594_n12342# 0.0023f
C914 a_n1500_n59307# a_n1500_n60543# 3.11f
C915 w_n1594_n11106# a_1500_n9770# 0.0023f
C916 a_1500_26074# w_n1594_27210# 0.0023f
C917 w_n1594_58110# a_1500_59446# 0.0023f
C918 a_1500_58210# w_n1594_58110# 0.0187f
C919 w_n1594_n61782# a_n1500_n63015# 0.0172f
C920 a_1500_43378# a_n1500_43281# 0.217f
C921 w_n1594_6198# a_n1558_5062# 0.0023f
C922 a_n1558_18658# w_n1594_18558# 0.0187f
C923 a_n1558_n29546# w_n1594_n29646# 0.0187f
C924 a_1500_38434# w_n1594_39570# 0.0023f
C925 a_n1500_51933# a_1500_52030# 0.217f
C926 w_n1594_n19758# a_n1558_n20894# 0.0023f
C927 a_n1500_n14811# w_n1594_n14814# 1.65f
C928 w_n1594_n27174# a_n1500_n27171# 1.65f
C929 a_n1558_3826# w_n1594_3726# 0.0187f
C930 a_1500_n46850# w_n1594_n45714# 0.0023f
C931 a_1500_24838# w_n1594_25974# 0.0023f
C932 a_n1500_n23463# a_n1558_n23366# 0.217f
C933 a_1500_n54266# w_n1594_n55602# 0.0023f
C934 w_n1594_n11106# a_1500_n12242# 0.0023f
C935 w_n1594_n13578# a_n1558_n12242# 0.0023f
C936 a_n1500_n14811# w_n1594_n16050# 0.0172f
C937 a_n1500_n63015# a_1500_n62918# 0.217f
C938 a_1500_33490# a_1500_34726# 0.0105f
C939 a_1500_n39434# a_1500_n40670# 0.0105f
C940 a_n1500_n40767# a_n1558_n40670# 0.217f
C941 w_n1594_60582# a_1500_61918# 0.0023f
C942 w_n1594_58110# a_n1558_59446# 0.0023f
C943 a_n1558_n45614# w_n1594_n44478# 0.0023f
C944 a_1500_22366# w_n1594_22266# 0.0187f
C945 w_n1594_n19758# a_n1558_n19658# 0.0187f
C946 a_n1500_58113# a_n1500_56877# 3.11f
C947 a_1500_58210# a_1500_56974# 0.0105f
C948 a_n1558_37198# a_n1558_35962# 0.0105f
C949 w_n1594_n58074# a_n1558_n56738# 0.0023f
C950 a_1500_n2354# w_n1594_n2454# 0.0187f
C951 a_1500_10006# w_n1594_8670# 0.0023f
C952 a_n1500_n32115# w_n1594_n33354# 0.0172f
C953 a_n1558_n33254# a_n1558_n34490# 0.0105f
C954 a_1500_40906# w_n1594_40806# 0.0187f
C955 w_n1594_16086# a_n1500_16089# 1.65f
C956 w_n1594_24738# a_n1558_26074# 0.0023f
C957 a_n1500_50697# w_n1594_50694# 1.65f
C958 a_1500_43378# a_1500_42142# 0.0105f
C959 a_n1558_n30782# w_n1594_n32118# 0.0023f
C960 a_n1558_n30782# w_n1594_n30882# 0.0187f
C961 a_1500_37198# w_n1594_38334# 0.0023f
C962 a_n1500_n23463# w_n1594_n22230# 0.0172f
C963 a_n1500_n24699# a_1500_n24602# 0.217f
C964 a_n1500_n6159# w_n1594_n4926# 0.0172f
C965 w_n1594_11142# a_1500_11242# 0.0187f
C966 a_n1558_1354# w_n1594_1254# 0.0187f
C967 w_n1594_8670# a_1500_7534# 0.0023f
C968 a_n1558_21130# a_n1558_22366# 0.0105f
C969 w_n1594_n43242# a_1500_n44378# 0.0023f
C970 a_n1500_n6159# a_n1500_n7395# 3.11f
C971 a_1500_n29546# a_1500_n28310# 0.0105f
C972 a_1500_n18422# a_n1500_n18519# 0.217f
C973 a_n1558_58210# a_n1558_59446# 0.0105f
C974 a_n1558_42142# w_n1594_43278# 0.0023f
C975 w_n1594_n40770# a_1500_n39434# 0.0023f
C976 w_n1594_n59310# a_n1558_n57974# 0.0023f
C977 a_n1500_n48183# a_1500_n48086# 0.217f
C978 a_n1500_n23463# w_n1594_n23466# 1.65f
C979 w_n1594_11142# a_1500_12478# 0.0023f
C980 a_n1558_n49322# w_n1594_n50658# 0.0023f
C981 w_n1594_37098# a_n1558_38434# 0.0023f
C982 a_1500_n17186# w_n1594_n16050# 0.0023f
C983 w_n1594_39570# a_n1558_39670# 0.0187f
C984 w_n1594_n38298# a_1500_n39434# 0.0023f
C985 a_n1500_22269# a_n1500_21033# 3.11f
C986 a_1500_31018# w_n1594_30918# 0.0187f
C987 a_n1558_n15950# a_n1500_n16047# 0.217f
C988 a_n1500_n51891# a_n1558_n51794# 0.217f
C989 a_1500_n50558# a_1500_n51794# 0.0105f
C990 a_1500_n29546# w_n1594_n28410# 0.0023f
C991 a_1500_n18422# w_n1594_n17286# 0.0023f
C992 a_n1500_35865# a_1500_35962# 0.217f
C993 a_n1558_43378# a_n1558_42142# 0.0105f
C994 w_n1594_61818# a_1500_60682# 0.0023f
C995 w_n1594_18# a_1500_n1118# 0.0023f
C996 a_n1500_60585# a_1500_60682# 0.217f
C997 w_n1594_48222# a_n1500_49461# 0.0172f
C998 a_n1500_n14811# a_n1500_n13575# 3.11f
C999 a_1500_11242# a_n1500_11145# 0.217f
C1000 w_n1594_1254# a_n1558_2590# 0.0023f
C1001 w_n1594_n43242# a_1500_n43142# 0.0187f
C1002 a_1500_53266# w_n1594_51930# 0.0023f
C1003 a_n1500_7437# a_n1500_8673# 3.11f
C1004 a_n1500_16089# a_n1500_17325# 3.11f
C1005 a_n1558_n9770# w_n1594_n8634# 0.0023f
C1006 w_n1594_n61782# a_n1500_n61779# 1.65f
C1007 a_n1500_n20991# a_n1558_n20894# 0.217f
C1008 w_n1594_n22230# a_n1500_n20991# 0.0172f
C1009 w_n1594_n55602# a_1500_n56738# 0.0023f
C1010 w_n1594_n25938# a_1500_n25838# 0.0187f
C1011 w_n1594_n1218# a_1500_118# 0.0023f
C1012 w_n1594_n27174# a_n1500_n25935# 0.0172f
C1013 a_n1558_23602# w_n1594_22266# 0.0023f
C1014 a_1500_n25838# w_n1594_n24702# 0.0023f
C1015 a_1500_n45614# w_n1594_n45714# 0.0187f
C1016 a_1500_n7298# a_n1500_n7395# 0.217f
C1017 w_n1594_59346# a_1500_60682# 0.0023f
C1018 a_n1500_25977# w_n1594_25974# 1.65f
C1019 w_n1594_n22230# a_1500_n20894# 0.0023f
C1020 a_1500_n50558# w_n1594_n49422# 0.0023f
C1021 a_n1558_22366# w_n1594_21030# 0.0023f
C1022 a_n1558_n61682# a_n1558_n62918# 0.0105f
C1023 a_1500_31018# w_n1594_32154# 0.0023f
C1024 a_n1558_n44378# w_n1594_n44478# 0.0187f
C1025 a_n1500_48225# a_n1500_46989# 3.11f
C1026 w_n1594_7434# a_1500_7534# 0.0187f
C1027 a_n1558_n27074# a_n1500_n27171# 0.217f
C1028 w_n1594_n17286# a_n1500_n16047# 0.0172f
C1029 a_1500_n27074# a_1500_n25838# 0.0105f
C1030 a_1500_43378# w_n1594_43278# 0.0187f
C1031 w_n1594_n56838# a_1500_n57974# 0.0023f
C1032 w_n1594_n60546# a_n1500_n61779# 0.0172f
C1033 w_n1594_23502# a_1500_24838# 0.0023f
C1034 a_n1500_n33351# a_1500_n33254# 0.217f
C1035 a_1500_22366# a_1500_23602# 0.0105f
C1036 a_n1500_22269# w_n1594_23502# 0.0172f
C1037 w_n1594_17322# a_1500_16186# 0.0023f
C1038 w_n1594_n34590# a_n1500_n35823# 0.0172f
C1039 a_n1500_4965# w_n1594_6198# 0.0172f
C1040 w_n1594_39570# a_n1500_40809# 0.0172f
C1041 a_n1558_37198# a_n1558_38434# 0.0105f
C1042 a_n1500_n43239# a_n1500_n44475# 3.11f
C1043 a_n1558_n29546# w_n1594_n30882# 0.0023f
C1044 a_n1500_43281# w_n1594_43278# 1.65f
C1045 a_1500_53266# w_n1594_54402# 0.0023f
C1046 w_n1594_60582# a_n1500_60585# 1.65f
C1047 a_n1558_13714# w_n1594_12378# 0.0023f
C1048 a_n1500_n32115# a_n1558_n32018# 0.217f
C1049 a_n1500_1257# w_n1594_1254# 1.65f
C1050 a_1500_n30782# a_1500_n32018# 0.0105f
C1051 a_1500_22366# w_n1594_21030# 0.0023f
C1052 a_1500_58210# a_1500_59446# 0.0105f
C1053 a_n1500_56877# a_n1500_55641# 3.11f
C1054 a_n1500_n37059# a_n1558_n36962# 0.217f
C1055 a_n1500_n11103# a_n1558_n11006# 0.217f
C1056 a_n1558_n46850# a_n1558_n48086# 0.0105f
C1057 w_n1594_n11106# a_n1558_n11006# 0.0187f
C1058 w_n1594_n38298# a_1500_n38198# 0.0187f
C1059 a_n1500_43281# a_n1500_44517# 3.11f
C1060 a_1500_1354# w_n1594_2490# 0.0023f
C1061 a_n1500_n7395# w_n1594_n7398# 1.65f
C1062 w_n1594_n44478# a_n1558_n43142# 0.0023f
C1063 a_n1558_45850# a_n1558_47086# 0.0105f
C1064 a_1500_13714# w_n1594_13614# 0.0187f
C1065 a_n1500_43281# a_n1558_43378# 0.217f
C1066 w_n1594_46986# a_n1500_45753# 0.0172f
C1067 a_1500_42142# w_n1594_43278# 0.0023f
C1068 w_n1594_n1218# a_n1558_118# 0.0023f
C1069 a_n1500_n17283# a_n1558_n17186# 0.217f
C1070 w_n1594_6198# a_1500_5062# 0.0023f
C1071 w_n1594_11142# a_n1500_11145# 1.65f
C1072 a_n1500_n4923# a_n1558_n4826# 0.217f
C1073 a_1500_n24602# w_n1594_n25938# 0.0023f
C1074 w_n1594_4962# a_1500_6298# 0.0023f
C1075 a_1500_n24602# w_n1594_n24702# 0.0187f
C1076 a_n1500_n58071# a_n1500_n59307# 3.11f
C1077 a_n1500_n14811# a_1500_n14714# 0.217f
C1078 w_n1594_4962# a_n1500_6201# 0.0172f
C1079 a_n1500_56877# a_n1558_56974# 0.217f
C1080 w_n1594_n42006# a_1500_n43142# 0.0023f
C1081 w_n1594_n43242# a_1500_n41906# 0.0023f
C1082 w_n1594_n61782# a_n1500_n60543# 0.0172f
C1083 a_n1500_n54363# a_n1500_n55599# 3.11f
C1084 w_n1594_n55602# a_1500_n55502# 0.0187f
C1085 a_n1500_39573# w_n1594_39570# 1.65f
C1086 w_n1594_33390# a_1500_34726# 0.0023f
C1087 w_n1594_n37062# a_n1500_n37059# 1.65f
C1088 a_1500_n44378# w_n1594_n45714# 0.0023f
C1089 a_1500_44614# a_1500_43378# 0.0105f
C1090 a_1500_n49322# w_n1594_n49422# 0.0187f
C1091 a_n1558_32254# w_n1594_33390# 0.0023f
C1092 a_n1500_n61779# a_1500_n61682# 0.217f
C1093 a_1500_n54266# w_n1594_n53130# 0.0023f
C1094 w_n1594_n14814# a_n1500_n16047# 0.0172f
C1095 a_1500_n38198# a_1500_n39434# 0.0105f
C1096 a_n1500_n39531# a_n1558_n39434# 0.217f
C1097 a_1500_47086# a_n1500_46989# 0.217f
C1098 a_n1500_n8631# a_n1500_n7395# 3.11f
C1099 a_1500_13714# a_1500_12478# 0.0105f
C1100 a_n1500_53169# a_n1500_54405# 3.11f
C1101 w_n1594_n16050# a_n1500_n16047# 1.65f
C1102 w_n1594_n56838# a_1500_n56738# 0.0187f
C1103 a_n1558_n6062# w_n1594_n6162# 0.0187f
C1104 a_1500_n54266# w_n1594_n54366# 0.0187f
C1105 a_n1500_n6159# w_n1594_n7398# 0.0172f
C1106 a_n1500_n11103# a_n1500_n9867# 3.11f
C1107 w_n1594_n60546# a_n1500_n60543# 1.65f
C1108 a_n1558_26074# w_n1594_25974# 0.0187f
C1109 a_1500_27310# w_n1594_27210# 0.0187f
C1110 w_n1594_n29646# a_n1500_n28407# 0.0172f
C1111 a_n1500_2493# a_n1558_2590# 0.217f
C1112 a_n1500_50697# w_n1594_49458# 0.0172f
C1113 w_n1594_n34590# a_n1500_n34587# 1.65f
C1114 a_n1558_12478# w_n1594_13614# 0.0023f
C1115 w_n1594_n12342# a_1500_n13478# 0.0023f
C1116 a_n1500_24741# a_n1558_24838# 0.217f
C1117 w_n1594_n11106# a_n1500_n9867# 0.0172f
C1118 w_n1594_n33354# a_n1500_n34587# 0.0172f
C1119 a_n1500_4965# a_n1558_5062# 0.217f
C1120 w_n1594_n35826# a_n1500_n37059# 0.0172f
C1121 w_n1594_n32118# a_n1558_n33254# 0.0023f
C1122 a_n1500_6201# a_n1500_7437# 3.11f
C1123 a_1500_13714# w_n1594_14850# 0.0023f
C1124 a_n1558_1354# a_n1558_118# 0.0105f
C1125 a_n1500_35865# w_n1594_34626# 0.0172f
C1126 w_n1594_6198# a_1500_7534# 0.0023f
C1127 a_1500_38434# w_n1594_38334# 0.0187f
C1128 a_1500_8770# a_n1500_8673# 0.217f
C1129 w_n1594_n27174# a_1500_n28310# 0.0023f
C1130 a_n1500_n46947# a_1500_n46850# 0.217f
C1131 w_n1594_24738# a_n1558_24838# 0.0187f
C1132 a_1500_49558# a_n1500_49461# 0.217f
C1133 w_n1594_n38298# a_1500_n36962# 0.0023f
C1134 w_n1594_17322# a_n1500_17325# 1.65f
C1135 w_n1594_n18522# a_1500_n17186# 0.0023f
C1136 a_1500_14950# w_n1594_13614# 0.0023f
C1137 a_n1558_n22130# a_n1500_n22227# 0.217f
C1138 a_n1500_33393# a_n1500_32157# 3.11f
C1139 a_1500_n23366# a_1500_n22130# 0.0105f
C1140 w_n1594_32154# a_n1558_33490# 0.0023f
C1141 a_n1500_1257# a_n1500_2493# 3.11f
C1142 a_n1500_n50655# a_n1558_n50558# 0.217f
C1143 a_1500_n49322# a_1500_n50558# 0.0105f
C1144 a_n1558_18658# a_n1558_17422# 0.0105f
C1145 a_1500_29782# w_n1594_30918# 0.0023f
C1146 a_1500_19894# a_n1500_19797# 0.217f
C1147 a_n1500_37101# a_n1500_35865# 3.11f
C1148 a_n1558_34726# w_n1594_35862# 0.0023f
C1149 a_n1500_58113# w_n1594_59346# 0.0172f
C1150 w_n1594_n1218# a_1500_n1118# 0.0187f
C1151 a_1500_n7298# w_n1594_n7398# 0.0187f
C1152 a_1500_n23366# w_n1594_n24702# 0.0023f
C1153 a_n1500_44517# w_n1594_43278# 0.0172f
C1154 a_n1500_39573# a_n1558_39670# 0.217f
C1155 a_n1500_n55599# a_n1500_n56835# 3.11f
C1156 w_n1594_45750# a_1500_47086# 0.0023f
C1157 w_n1594_n42006# a_1500_n41906# 0.0187f
C1158 a_1500_n6062# a_1500_n4826# 0.0105f
C1159 a_n1558_n15950# a_n1558_n17186# 0.0105f
C1160 a_1500_n18422# a_1500_n19658# 0.0105f
C1161 a_n1558_49558# a_n1500_49461# 0.217f
C1162 a_n1558_43378# w_n1594_43278# 0.0187f
C1163 w_n1594_n28410# a_n1558_n28310# 0.0187f
C1164 a_n1558_53266# a_n1558_54502# 0.0105f
C1165 w_n1594_48222# a_n1558_48322# 0.0187f
C1166 w_n1594_56874# a_1500_55738# 0.0023f
C1167 w_n1594_n37062# a_n1500_n35823# 0.0172f
C1168 a_1500_3826# a_1500_2590# 0.0105f
C1169 a_1500_42142# a_1500_40906# 0.0105f
C1170 a_n1500_n14811# a_n1558_n14714# 0.217f
C1171 a_1500_n48086# w_n1594_n49422# 0.0023f
C1172 w_n1594_12378# a_n1558_11242# 0.0023f
C1173 w_n1594_32154# a_n1500_33393# 0.0172f
C1174 w_n1594_38334# a_n1558_39670# 0.0023f
C1175 a_1500_n53030# w_n1594_n53130# 0.0187f
C1176 w_n1594_61818# a_n1558_60682# 0.0023f
C1177 a_n1558_n60446# a_n1558_n61682# 0.0105f
C1178 w_n1594_50694# a_n1558_50794# 0.0187f
C1179 w_n1594_11142# a_n1500_9909# 0.0172f
C1180 w_n1594_46986# a_n1558_45850# 0.0023f
C1181 a_n1558_n4826# w_n1594_n6162# 0.0023f
C1182 a_n1500_60585# a_n1558_60682# 0.217f
C1183 a_n1500_25977# a_n1558_26074# 0.217f
C1184 a_n1558_n3590# a_n1500_n3687# 0.217f
C1185 a_n1500_6201# a_n1558_6298# 0.217f
C1186 w_n1594_n63018# a_n1558_n62918# 0.0187f
C1187 a_n1500_n12339# a_1500_n12242# 0.217f
C1188 w_n1594_n56838# a_1500_n55502# 0.0023f
C1189 a_1500_n53030# w_n1594_n54366# 0.0023f
C1190 w_n1594_48222# a_1500_48322# 0.0187f
C1191 w_n1594_n60546# a_n1500_n59307# 0.0172f
C1192 a_n1500_n48183# w_n1594_n46950# 0.0172f
C1193 a_1500_14950# w_n1594_14850# 0.0187f
C1194 w_n1594_n34590# a_n1500_n33351# 0.0172f
C1195 a_n1500_29685# w_n1594_28446# 0.0172f
C1196 w_n1594_n33354# a_n1500_n33351# 1.65f
C1197 w_n1594_59346# a_n1558_60682# 0.0023f
C1198 a_n1500_n42003# a_n1500_n43239# 3.11f
C1199 w_n1594_n37062# a_n1500_n38295# 0.0172f
C1200 w_n1594_n35826# a_n1500_n35823# 1.65f
C1201 w_n1594_n19758# a_n1558_n18422# 0.0023f
C1202 a_n1500_n30879# a_n1558_n30782# 0.217f
C1203 a_1500_n29546# a_1500_n30782# 0.0105f
C1204 a_n1500_40809# w_n1594_42042# 0.0172f
C1205 a_n1500_n11103# w_n1594_n12342# 0.0172f
C1206 w_n1594_n2454# a_n1558_n1118# 0.0023f
C1207 a_n1500_27213# w_n1594_27210# 1.65f
C1208 a_n1558_n8534# w_n1594_n7398# 0.0023f
C1209 a_1500_44614# w_n1594_43278# 0.0023f
C1210 a_1500_n32018# a_1500_n33254# 0.0105f
C1211 w_n1594_n17286# a_n1558_n17186# 0.0187f
C1212 a_n1558_33490# w_n1594_34626# 0.0023f
C1213 a_n1500_37101# w_n1594_38334# 0.0172f
C1214 a_n1500_n35823# a_n1558_n35726# 0.217f
C1215 w_n1594_18# a_n1500_21# 1.65f
C1216 a_1500_n34490# a_1500_n35726# 0.0105f
C1217 a_n1500_n49419# w_n1594_n48186# 0.0172f
C1218 w_n1594_n27174# a_1500_n27074# 0.0187f
C1219 a_n1558_n45614# a_n1558_n46850# 0.0105f
C1220 a_n1558_12478# w_n1594_11142# 0.0023f
C1221 w_n1594_n13578# a_1500_n13478# 0.0187f
C1222 a_n1500_39573# a_n1500_40809# 3.11f
C1223 w_n1594_39570# a_n1500_38337# 0.0172f
C1224 a_1500_n8534# w_n1594_n8634# 0.0187f
C1225 a_n1500_n53127# w_n1594_n51894# 0.0172f
C1226 w_n1594_n17286# a_1500_n15950# 0.0023f
C1227 w_n1594_30918# a_n1558_29782# 0.0023f
C1228 a_n1500_n4923# a_1500_n4826# 0.217f
C1229 a_n1500_11145# a_n1500_9909# 3.11f
C1230 w_n1594_28446# a_n1558_28546# 0.0187f
C1231 a_1500_44614# a_n1500_44517# 0.217f
C1232 w_n1594_12378# a_n1500_13617# 0.0172f
C1233 a_n1558_7534# w_n1594_8670# 0.0023f
C1234 a_1500_n35726# a_1500_n36962# 0.0105f
C1235 a_n1500_33393# w_n1594_34626# 0.0172f
C1236 a_n1500_n24699# w_n1594_n23466# 0.0172f
C1237 w_n1594_28446# a_1500_28546# 0.0187f
C1238 w_n1594_n39534# a_n1500_n40767# 0.0172f
C1239 a_n1558_55738# w_n1594_54402# 0.0023f
C1240 w_n1594_n20994# a_n1558_n22130# 0.0023f
C1241 w_n1594_n18522# a_1500_n18422# 0.0187f
C1242 a_n1500_n56835# a_n1500_n58071# 3.11f
C1243 a_1500_38434# a_n1500_38337# 0.217f
C1244 a_n1558_n8534# a_n1500_n8631# 0.217f
C1245 w_n1594_56874# a_1500_56974# 0.0187f
C1246 a_n1500_16089# a_n1500_14853# 3.11f
C1247 a_n1558_58210# w_n1594_56874# 0.0023f
C1248 w_n1594_n42006# a_1500_n40670# 0.0023f
C1249 a_n1500_n53127# a_n1500_n54363# 3.11f
C1250 a_n1558_55738# w_n1594_55638# 0.0187f
C1251 w_n1594_n28410# a_n1558_n27074# 0.0023f
C1252 a_n1500_34629# w_n1594_33390# 0.0172f
C1253 a_n1500_n8631# w_n1594_n7398# 0.0172f
C1254 a_n1558_n2354# a_n1500_n2451# 0.217f
C1255 w_n1594_n22230# a_n1500_n22227# 1.65f
C1256 a_1500_54502# w_n1594_54402# 0.0187f
C1257 a_n1558_n9770# w_n1594_n11106# 0.0023f
C1258 a_1500_50794# w_n1594_51930# 0.0023f
C1259 a_1500_1354# w_n1594_18# 0.0023f
C1260 a_1500_n51794# w_n1594_n53130# 0.0023f
C1261 a_n1500_n60543# a_1500_n60446# 0.217f
C1262 a_1500_n36962# a_1500_n38198# 0.0105f
C1263 a_n1500_n38295# a_n1558_n38198# 0.217f
C1264 a_n1500_60585# a_n1500_59349# 3.11f
C1265 a_1500_61918# a_n1500_61821# 0.217f
C1266 a_1500_54502# w_n1594_55638# 0.0023f
C1267 w_n1594_n63018# a_n1558_n61682# 0.0023f
C1268 a_n1500_4965# a_1500_5062# 0.217f
C1269 a_n1500_34629# a_n1558_34726# 0.217f
C1270 w_n1594_n54366# a_1500_n55502# 0.0023f
C1271 a_n1500_n22227# w_n1594_n23466# 0.0172f
C1272 a_n1558_19894# a_n1500_19797# 0.217f
C1273 a_1500_19894# w_n1594_21030# 0.0023f
C1274 w_n1594_n1218# a_n1500_n2451# 0.0172f
C1275 a_1500_53266# a_n1500_53169# 0.217f
C1276 a_n1500_n46947# w_n1594_n46950# 1.65f
C1277 w_n1594_59346# a_n1500_59349# 1.65f
C1278 a_n1500_27213# a_n1558_27310# 0.217f
C1279 w_n1594_n35826# a_n1500_n34587# 0.0172f
C1280 a_n1500_18561# a_n1558_18658# 0.217f
C1281 a_n1558_32254# a_n1558_31018# 0.0105f
C1282 a_1500_31018# a_1500_29782# 0.0105f
C1283 w_n1594_n16050# a_n1558_n17186# 0.0023f
C1284 a_1500_53266# a_1500_52030# 0.0105f
C1285 a_n1500_27213# a_n1500_28449# 3.11f
C1286 a_n1558_21130# w_n1594_22266# 0.0023f
C1287 a_n1500_39573# w_n1594_38334# 0.0172f
C1288 w_n1594_n58074# a_n1500_n59307# 0.0172f
C1289 a_1500_39670# a_1500_40906# 0.0105f
C1290 w_n1594_n25938# a_n1558_n27074# 0.0023f
C1291 a_n1500_n45711# a_1500_n45614# 0.217f
C1292 a_n1500_n48183# w_n1594_n48186# 1.65f
C1293 a_n1558_24838# w_n1594_25974# 0.0023f
C1294 a_n1558_7534# w_n1594_7434# 0.0187f
C1295 a_1500_n15950# w_n1594_n14814# 0.0023f
C1296 a_n1500_17325# w_n1594_18558# 0.0172f
C1297 a_n1500_n51891# w_n1594_n51894# 1.65f
C1298 w_n1594_n16050# a_1500_n15950# 0.0187f
C1299 a_n1558_n8534# w_n1594_n9870# 0.0023f
C1300 w_n1594_n40770# a_n1558_n41906# 0.0023f
C1301 a_n1500_16089# a_n1558_16186# 0.217f
C1302 w_n1594_n59310# a_n1500_n60543# 0.0172f
C1303 a_n1500_51933# w_n1594_53166# 0.0172f
C1304 a_1500_n48086# a_1500_n49322# 0.0105f
C1305 a_n1500_n49419# a_n1558_n49322# 0.217f
C1306 a_1500_n24602# a_1500_n25838# 0.0105f
C1307 a_n1500_n51891# w_n1594_n50658# 0.0172f
C1308 a_n1500_n7395# a_n1558_n7298# 0.217f
C1309 w_n1594_3726# a_n1500_2493# 0.0172f
C1310 a_n1500_12381# w_n1594_12378# 1.65f
C1311 a_n1500_8673# a_n1500_9909# 3.11f
C1312 a_n1558_n23366# w_n1594_n24702# 0.0023f
C1313 w_n1594_n39534# a_n1500_n39531# 1.65f
C1314 a_n1558_n19658# a_n1500_n19755# 0.217f
C1315 a_n1500_37101# a_n1500_38337# 3.11f
C1316 a_n1500_n25935# a_n1558_n25838# 0.217f
C1317 a_n1500_14853# a_n1500_13617# 3.11f
C1318 a_n1500_7437# w_n1594_8670# 0.0172f
C1319 a_1500_48322# a_1500_49558# 0.0105f
C1320 a_n1500_50697# a_n1558_50794# 0.217f
C1321 w_n1594_21030# a_n1500_19797# 0.0172f
C1322 a_n1500_29685# w_n1594_29682# 1.65f
C1323 a_1500_n4826# w_n1594_n6162# 0.0023f
C1324 a_n1558_21130# a_n1558_19894# 0.0105f
C1325 w_n1594_n22230# a_1500_n22130# 0.0187f
C1326 a_n1558_n3590# w_n1594_n2454# 0.0023f
C1327 w_n1594_16086# a_n1558_14950# 0.0023f
C1328 a_1500_23602# w_n1594_22266# 0.0023f
C1329 a_n1558_n59210# a_n1558_n60446# 0.0105f
C1330 a_n1558_48322# a_n1558_49558# 0.0105f
C1331 w_n1594_49458# a_n1558_50794# 0.0023f
C1332 a_n1500_23505# a_n1558_23602# 0.217f
C1333 a_n1558_13714# a_n1500_13617# 0.217f
C1334 a_1500_58210# w_n1594_56874# 0.0023f
C1335 a_1500_n22130# w_n1594_n23466# 0.0023f
C1336 w_n1594_n61782# a_1500_n62918# 0.0023f
C1337 a_n1558_n20894# w_n1594_n20994# 0.0187f
C1338 a_n1558_40906# w_n1594_39570# 0.0023f
C1339 a_n1500_n30879# w_n1594_n29646# 0.0172f
C1340 a_1500_54502# a_1500_55738# 0.0105f
C1341 a_n1500_n8631# w_n1594_n9870# 0.0172f
C1342 a_n1558_n55502# w_n1594_n55602# 0.0187f
C1343 a_n1500_n45711# w_n1594_n46950# 0.0172f
C1344 a_n1558_28546# w_n1594_29682# 0.0023f
C1345 w_n1594_61818# a_n1500_61821# 1.65f
C1346 w_n1594_11142# a_n1558_10006# 0.0023f
C1347 w_n1594_n4926# a_1500_n6062# 0.0023f
C1348 w_n1594_9906# a_1500_11242# 0.0023f
C1349 a_n1500_n40767# a_n1500_n42003# 3.11f
C1350 a_n1558_n19658# w_n1594_n20994# 0.0023f
C1351 a_n1500_n29643# a_n1558_n29546# 0.217f
C1352 a_n1500_60585# a_n1500_61821# 3.11f
C1353 a_n1558_52030# w_n1594_53166# 0.0023f
C1354 w_n1594_48222# a_1500_49558# 0.0023f
C1355 a_1500_28546# w_n1594_29682# 0.0023f
C1356 a_n1500_53169# w_n1594_53166# 1.65f
C1357 w_n1594_n58074# a_n1500_n58071# 1.65f
C1358 a_1500_n33254# a_1500_n34490# 0.0105f
C1359 a_n1500_n34587# a_n1558_n34490# 0.217f
C1360 w_n1594_n1218# a_n1500_21# 0.0172f
C1361 a_1500_n32018# w_n1594_n33354# 0.0023f
C1362 a_1500_14950# a_1500_13714# 0.0105f
C1363 a_n1558_n44378# a_n1558_n45614# 0.0105f
C1364 a_n1500_n46947# w_n1594_n48186# 0.0172f
C1365 a_n1500_n32115# w_n1594_n32118# 1.65f
C1366 a_n1500_n32115# w_n1594_n30882# 0.0172f
C1367 a_1500_21130# a_1500_22366# 0.0105f
C1368 a_n1500_n50655# w_n1594_n51894# 0.0172f
C1369 a_1500_52030# w_n1594_53166# 0.0023f
C1370 w_n1594_21030# a_n1558_19894# 0.0023f
C1371 a_1500_n4826# a_1500_n3590# 0.0105f
C1372 w_n1594_n40770# a_n1558_n40670# 0.0187f
C1373 a_n1558_21130# w_n1594_21030# 0.0187f
C1374 a_n1500_7437# w_n1594_7434# 1.65f
C1375 w_n1594_n59310# a_n1500_n59307# 1.65f
C1376 w_n1594_14850# a_1500_16186# 0.0023f
C1377 a_n1500_n50655# w_n1594_n50658# 1.65f
C1378 a_1500_8770# w_n1594_9906# 0.0023f
C1379 a_1500_27310# a_1500_26074# 0.0105f
C1380 w_n1594_n12342# a_n1500_n13575# 0.0172f
C1381 a_n1558_7534# w_n1594_6198# 0.0023f
C1382 a_n1558_24838# w_n1594_23502# 0.0023f
C1383 w_n1594_48222# a_n1558_49558# 0.0023f
C1384 w_n1594_29682# a_n1558_31018# 0.0023f
C1385 a_n1558_n13478# w_n1594_n14814# 0.0023f
C1386 w_n1594_n39534# a_n1500_n38295# 0.0172f
C1387 a_n1500_33393# a_n1558_33490# 0.217f
C1388 w_n1594_54402# a_n1558_54502# 0.0187f
C1389 a_n1500_39573# a_n1500_38337# 3.11f
C1390 a_n1558_n2354# w_n1594_n2454# 0.0187f
C1391 a_n1500_n51891# a_n1500_n53127# 3.11f
C1392 a_n1500_n6159# a_1500_n6062# 0.217f
C1393 a_1500_34726# w_n1594_35862# 0.0023f
C1394 a_n1558_35962# w_n1594_34626# 0.0023f
C1395 w_n1594_46986# a_n1558_47086# 0.0187f
C1396 w_n1594_1254# a_1500_118# 0.0023f
C1397 w_n1594_24738# a_n1558_23602# 0.0023f
C1398 a_1500_19894# a_1500_18658# 0.0105f
C1399 w_n1594_55638# a_n1558_54502# 0.0023f
C1400 w_n1594_1254# a_n1500_2493# 0.0172f
C1401 a_1500_n44378# a_n1500_n44475# 0.217f
C1402 a_n1500_n4923# w_n1594_n4926# 1.65f
C1403 w_n1594_38334# a_n1500_38337# 1.65f
C1404 a_n1500_n14811# a_n1500_n16047# 3.11f
C1405 a_n1500_n59307# a_1500_n59210# 0.217f
C1406 a_n1558_40906# a_n1558_39670# 0.0105f
C1407 a_n1500_n18519# a_n1558_n18422# 0.217f
C1408 a_1500_n18422# a_1500_n17186# 0.0105f
C1409 w_n1594_n61782# a_1500_n61682# 0.0187f
C1410 a_1500_45850# w_n1594_44514# 0.0023f
C1411 a_n1500_n29643# w_n1594_n29646# 1.65f
C1412 w_n1594_n27174# a_1500_n25838# 0.0023f
C1413 w_n1594_32154# a_1500_33490# 0.0023f
C1414 a_1500_n9770# w_n1594_n9870# 0.0187f
C1415 w_n1594_39570# a_n1558_38434# 0.0023f
C1416 a_n1558_n54266# w_n1594_n55602# 0.0023f
C1417 w_n1594_n11106# a_n1558_n12242# 0.0023f
C1418 a_n1558_n46850# w_n1594_n45714# 0.0023f
C1419 a_1500_n62918# VSUBS 0.638f
C1420 a_n1558_n62918# VSUBS 0.638f
C1421 a_n1500_n63015# VSUBS 5.03f
C1422 a_1500_n61682# VSUBS 0.625f
C1423 a_n1558_n61682# VSUBS 0.625f
C1424 a_n1500_n61779# VSUBS 3.31f
C1425 a_1500_n60446# VSUBS 0.625f
C1426 a_n1558_n60446# VSUBS 0.625f
C1427 a_n1500_n60543# VSUBS 3.31f
C1428 a_1500_n59210# VSUBS 0.625f
C1429 a_n1558_n59210# VSUBS 0.625f
C1430 a_n1500_n59307# VSUBS 3.31f
C1431 a_1500_n57974# VSUBS 0.625f
C1432 a_n1558_n57974# VSUBS 0.625f
C1433 a_n1500_n58071# VSUBS 3.31f
C1434 a_1500_n56738# VSUBS 0.625f
C1435 a_n1558_n56738# VSUBS 0.625f
C1436 a_n1500_n56835# VSUBS 3.31f
C1437 a_1500_n55502# VSUBS 0.625f
C1438 a_n1558_n55502# VSUBS 0.625f
C1439 a_n1500_n55599# VSUBS 3.31f
C1440 a_1500_n54266# VSUBS 0.625f
C1441 a_n1558_n54266# VSUBS 0.625f
C1442 a_n1500_n54363# VSUBS 3.31f
C1443 a_1500_n53030# VSUBS 0.625f
C1444 a_n1558_n53030# VSUBS 0.625f
C1445 a_n1500_n53127# VSUBS 3.31f
C1446 a_1500_n51794# VSUBS 0.625f
C1447 a_n1558_n51794# VSUBS 0.625f
C1448 a_n1500_n51891# VSUBS 3.31f
C1449 a_1500_n50558# VSUBS 0.625f
C1450 a_n1558_n50558# VSUBS 0.625f
C1451 a_n1500_n50655# VSUBS 3.31f
C1452 a_1500_n49322# VSUBS 0.625f
C1453 a_n1558_n49322# VSUBS 0.625f
C1454 a_n1500_n49419# VSUBS 3.31f
C1455 a_1500_n48086# VSUBS 0.625f
C1456 a_n1558_n48086# VSUBS 0.625f
C1457 a_n1500_n48183# VSUBS 3.31f
C1458 a_1500_n46850# VSUBS 0.625f
C1459 a_n1558_n46850# VSUBS 0.625f
C1460 a_n1500_n46947# VSUBS 3.31f
C1461 a_1500_n45614# VSUBS 0.625f
C1462 a_n1558_n45614# VSUBS 0.625f
C1463 a_n1500_n45711# VSUBS 3.31f
C1464 a_1500_n44378# VSUBS 0.625f
C1465 a_n1558_n44378# VSUBS 0.625f
C1466 a_n1500_n44475# VSUBS 3.31f
C1467 a_1500_n43142# VSUBS 0.625f
C1468 a_n1558_n43142# VSUBS 0.625f
C1469 a_n1500_n43239# VSUBS 3.31f
C1470 a_1500_n41906# VSUBS 0.625f
C1471 a_n1558_n41906# VSUBS 0.625f
C1472 a_n1500_n42003# VSUBS 3.31f
C1473 a_1500_n40670# VSUBS 0.625f
C1474 a_n1558_n40670# VSUBS 0.625f
C1475 a_n1500_n40767# VSUBS 3.31f
C1476 a_1500_n39434# VSUBS 0.625f
C1477 a_n1558_n39434# VSUBS 0.625f
C1478 a_n1500_n39531# VSUBS 3.31f
C1479 a_1500_n38198# VSUBS 0.625f
C1480 a_n1558_n38198# VSUBS 0.625f
C1481 a_n1500_n38295# VSUBS 3.31f
C1482 a_1500_n36962# VSUBS 0.625f
C1483 a_n1558_n36962# VSUBS 0.625f
C1484 a_n1500_n37059# VSUBS 3.31f
C1485 a_1500_n35726# VSUBS 0.625f
C1486 a_n1558_n35726# VSUBS 0.625f
C1487 a_n1500_n35823# VSUBS 3.31f
C1488 a_1500_n34490# VSUBS 0.625f
C1489 a_n1558_n34490# VSUBS 0.625f
C1490 a_n1500_n34587# VSUBS 3.31f
C1491 a_1500_n33254# VSUBS 0.625f
C1492 a_n1558_n33254# VSUBS 0.625f
C1493 a_n1500_n33351# VSUBS 3.31f
C1494 a_1500_n32018# VSUBS 0.625f
C1495 a_n1558_n32018# VSUBS 0.625f
C1496 a_n1500_n32115# VSUBS 3.31f
C1497 a_1500_n30782# VSUBS 0.625f
C1498 a_n1558_n30782# VSUBS 0.625f
C1499 a_n1500_n30879# VSUBS 3.31f
C1500 a_1500_n29546# VSUBS 0.625f
C1501 a_n1558_n29546# VSUBS 0.625f
C1502 a_n1500_n29643# VSUBS 3.31f
C1503 a_1500_n28310# VSUBS 0.625f
C1504 a_n1558_n28310# VSUBS 0.625f
C1505 a_n1500_n28407# VSUBS 3.31f
C1506 a_1500_n27074# VSUBS 0.625f
C1507 a_n1558_n27074# VSUBS 0.625f
C1508 a_n1500_n27171# VSUBS 3.31f
C1509 a_1500_n25838# VSUBS 0.625f
C1510 a_n1558_n25838# VSUBS 0.625f
C1511 a_n1500_n25935# VSUBS 3.31f
C1512 a_1500_n24602# VSUBS 0.625f
C1513 a_n1558_n24602# VSUBS 0.625f
C1514 a_n1500_n24699# VSUBS 3.31f
C1515 a_1500_n23366# VSUBS 0.625f
C1516 a_n1558_n23366# VSUBS 0.625f
C1517 a_n1500_n23463# VSUBS 3.31f
C1518 a_1500_n22130# VSUBS 0.625f
C1519 a_n1558_n22130# VSUBS 0.625f
C1520 a_n1500_n22227# VSUBS 3.31f
C1521 a_1500_n20894# VSUBS 0.625f
C1522 a_n1558_n20894# VSUBS 0.625f
C1523 a_n1500_n20991# VSUBS 3.31f
C1524 a_1500_n19658# VSUBS 0.625f
C1525 a_n1558_n19658# VSUBS 0.625f
C1526 a_n1500_n19755# VSUBS 3.31f
C1527 a_1500_n18422# VSUBS 0.625f
C1528 a_n1558_n18422# VSUBS 0.625f
C1529 a_n1500_n18519# VSUBS 3.31f
C1530 a_1500_n17186# VSUBS 0.625f
C1531 a_n1558_n17186# VSUBS 0.625f
C1532 a_n1500_n17283# VSUBS 3.31f
C1533 a_1500_n15950# VSUBS 0.625f
C1534 a_n1558_n15950# VSUBS 0.625f
C1535 a_n1500_n16047# VSUBS 3.31f
C1536 a_1500_n14714# VSUBS 0.625f
C1537 a_n1558_n14714# VSUBS 0.625f
C1538 a_n1500_n14811# VSUBS 3.31f
C1539 a_1500_n13478# VSUBS 0.625f
C1540 a_n1558_n13478# VSUBS 0.625f
C1541 a_n1500_n13575# VSUBS 3.31f
C1542 a_1500_n12242# VSUBS 0.625f
C1543 a_n1558_n12242# VSUBS 0.625f
C1544 a_n1500_n12339# VSUBS 3.31f
C1545 a_1500_n11006# VSUBS 0.625f
C1546 a_n1558_n11006# VSUBS 0.625f
C1547 a_n1500_n11103# VSUBS 3.31f
C1548 a_1500_n9770# VSUBS 0.625f
C1549 a_n1558_n9770# VSUBS 0.625f
C1550 a_n1500_n9867# VSUBS 3.31f
C1551 a_1500_n8534# VSUBS 0.625f
C1552 a_n1558_n8534# VSUBS 0.625f
C1553 a_n1500_n8631# VSUBS 3.31f
C1554 a_1500_n7298# VSUBS 0.625f
C1555 a_n1558_n7298# VSUBS 0.625f
C1556 a_n1500_n7395# VSUBS 3.31f
C1557 a_1500_n6062# VSUBS 0.625f
C1558 a_n1558_n6062# VSUBS 0.625f
C1559 a_n1500_n6159# VSUBS 3.31f
C1560 a_1500_n4826# VSUBS 0.625f
C1561 a_n1558_n4826# VSUBS 0.625f
C1562 a_n1500_n4923# VSUBS 3.31f
C1563 a_1500_n3590# VSUBS 0.625f
C1564 a_n1558_n3590# VSUBS 0.625f
C1565 a_n1500_n3687# VSUBS 3.31f
C1566 a_1500_n2354# VSUBS 0.625f
C1567 a_n1558_n2354# VSUBS 0.625f
C1568 a_n1500_n2451# VSUBS 3.31f
C1569 a_1500_n1118# VSUBS 0.625f
C1570 a_n1558_n1118# VSUBS 0.625f
C1571 a_n1500_n1215# VSUBS 3.31f
C1572 a_1500_118# VSUBS 0.625f
C1573 a_n1558_118# VSUBS 0.625f
C1574 a_n1500_21# VSUBS 3.31f
C1575 a_1500_1354# VSUBS 0.625f
C1576 a_n1558_1354# VSUBS 0.625f
C1577 a_n1500_1257# VSUBS 3.31f
C1578 a_1500_2590# VSUBS 0.625f
C1579 a_n1558_2590# VSUBS 0.625f
C1580 a_n1500_2493# VSUBS 3.31f
C1581 a_1500_3826# VSUBS 0.625f
C1582 a_n1558_3826# VSUBS 0.625f
C1583 a_n1500_3729# VSUBS 3.31f
C1584 a_1500_5062# VSUBS 0.625f
C1585 a_n1558_5062# VSUBS 0.625f
C1586 a_n1500_4965# VSUBS 3.31f
C1587 a_1500_6298# VSUBS 0.625f
C1588 a_n1558_6298# VSUBS 0.625f
C1589 a_n1500_6201# VSUBS 3.31f
C1590 a_1500_7534# VSUBS 0.625f
C1591 a_n1558_7534# VSUBS 0.625f
C1592 a_n1500_7437# VSUBS 3.31f
C1593 a_1500_8770# VSUBS 0.625f
C1594 a_n1558_8770# VSUBS 0.625f
C1595 a_n1500_8673# VSUBS 3.31f
C1596 a_1500_10006# VSUBS 0.625f
C1597 a_n1558_10006# VSUBS 0.625f
C1598 a_n1500_9909# VSUBS 3.31f
C1599 a_1500_11242# VSUBS 0.625f
C1600 a_n1558_11242# VSUBS 0.625f
C1601 a_n1500_11145# VSUBS 3.31f
C1602 a_1500_12478# VSUBS 0.625f
C1603 a_n1558_12478# VSUBS 0.625f
C1604 a_n1500_12381# VSUBS 3.31f
C1605 a_1500_13714# VSUBS 0.625f
C1606 a_n1558_13714# VSUBS 0.625f
C1607 a_n1500_13617# VSUBS 3.31f
C1608 a_1500_14950# VSUBS 0.625f
C1609 a_n1558_14950# VSUBS 0.625f
C1610 a_n1500_14853# VSUBS 3.31f
C1611 a_1500_16186# VSUBS 0.625f
C1612 a_n1558_16186# VSUBS 0.625f
C1613 a_n1500_16089# VSUBS 3.31f
C1614 a_1500_17422# VSUBS 0.625f
C1615 a_n1558_17422# VSUBS 0.625f
C1616 a_n1500_17325# VSUBS 3.31f
C1617 a_1500_18658# VSUBS 0.625f
C1618 a_n1558_18658# VSUBS 0.625f
C1619 a_n1500_18561# VSUBS 3.31f
C1620 a_1500_19894# VSUBS 0.625f
C1621 a_n1558_19894# VSUBS 0.625f
C1622 a_n1500_19797# VSUBS 3.31f
C1623 a_1500_21130# VSUBS 0.625f
C1624 a_n1558_21130# VSUBS 0.625f
C1625 a_n1500_21033# VSUBS 3.31f
C1626 a_1500_22366# VSUBS 0.625f
C1627 a_n1558_22366# VSUBS 0.625f
C1628 a_n1500_22269# VSUBS 3.31f
C1629 a_1500_23602# VSUBS 0.625f
C1630 a_n1558_23602# VSUBS 0.625f
C1631 a_n1500_23505# VSUBS 3.31f
C1632 a_1500_24838# VSUBS 0.625f
C1633 a_n1558_24838# VSUBS 0.625f
C1634 a_n1500_24741# VSUBS 3.31f
C1635 a_1500_26074# VSUBS 0.625f
C1636 a_n1558_26074# VSUBS 0.625f
C1637 a_n1500_25977# VSUBS 3.31f
C1638 a_1500_27310# VSUBS 0.625f
C1639 a_n1558_27310# VSUBS 0.625f
C1640 a_n1500_27213# VSUBS 3.31f
C1641 a_1500_28546# VSUBS 0.625f
C1642 a_n1558_28546# VSUBS 0.625f
C1643 a_n1500_28449# VSUBS 3.31f
C1644 a_1500_29782# VSUBS 0.625f
C1645 a_n1558_29782# VSUBS 0.625f
C1646 a_n1500_29685# VSUBS 3.31f
C1647 a_1500_31018# VSUBS 0.625f
C1648 a_n1558_31018# VSUBS 0.625f
C1649 a_n1500_30921# VSUBS 3.31f
C1650 a_1500_32254# VSUBS 0.625f
C1651 a_n1558_32254# VSUBS 0.625f
C1652 a_n1500_32157# VSUBS 3.31f
C1653 a_1500_33490# VSUBS 0.625f
C1654 a_n1558_33490# VSUBS 0.625f
C1655 a_n1500_33393# VSUBS 3.31f
C1656 a_1500_34726# VSUBS 0.625f
C1657 a_n1558_34726# VSUBS 0.625f
C1658 a_n1500_34629# VSUBS 3.31f
C1659 a_1500_35962# VSUBS 0.625f
C1660 a_n1558_35962# VSUBS 0.625f
C1661 a_n1500_35865# VSUBS 3.31f
C1662 a_1500_37198# VSUBS 0.625f
C1663 a_n1558_37198# VSUBS 0.625f
C1664 a_n1500_37101# VSUBS 3.31f
C1665 a_1500_38434# VSUBS 0.625f
C1666 a_n1558_38434# VSUBS 0.625f
C1667 a_n1500_38337# VSUBS 3.31f
C1668 a_1500_39670# VSUBS 0.625f
C1669 a_n1558_39670# VSUBS 0.625f
C1670 a_n1500_39573# VSUBS 3.31f
C1671 a_1500_40906# VSUBS 0.625f
C1672 a_n1558_40906# VSUBS 0.625f
C1673 a_n1500_40809# VSUBS 3.31f
C1674 a_1500_42142# VSUBS 0.625f
C1675 a_n1558_42142# VSUBS 0.625f
C1676 a_n1500_42045# VSUBS 3.31f
C1677 a_1500_43378# VSUBS 0.625f
C1678 a_n1558_43378# VSUBS 0.625f
C1679 a_n1500_43281# VSUBS 3.31f
C1680 a_1500_44614# VSUBS 0.625f
C1681 a_n1558_44614# VSUBS 0.625f
C1682 a_n1500_44517# VSUBS 3.31f
C1683 a_1500_45850# VSUBS 0.625f
C1684 a_n1558_45850# VSUBS 0.625f
C1685 a_n1500_45753# VSUBS 3.31f
C1686 a_1500_47086# VSUBS 0.625f
C1687 a_n1558_47086# VSUBS 0.625f
C1688 a_n1500_46989# VSUBS 3.31f
C1689 a_1500_48322# VSUBS 0.625f
C1690 a_n1558_48322# VSUBS 0.625f
C1691 a_n1500_48225# VSUBS 3.31f
C1692 a_1500_49558# VSUBS 0.625f
C1693 a_n1558_49558# VSUBS 0.625f
C1694 a_n1500_49461# VSUBS 3.31f
C1695 a_1500_50794# VSUBS 0.625f
C1696 a_n1558_50794# VSUBS 0.625f
C1697 a_n1500_50697# VSUBS 3.31f
C1698 a_1500_52030# VSUBS 0.625f
C1699 a_n1558_52030# VSUBS 0.625f
C1700 a_n1500_51933# VSUBS 3.31f
C1701 a_1500_53266# VSUBS 0.625f
C1702 a_n1558_53266# VSUBS 0.625f
C1703 a_n1500_53169# VSUBS 3.31f
C1704 a_1500_54502# VSUBS 0.625f
C1705 a_n1558_54502# VSUBS 0.625f
C1706 a_n1500_54405# VSUBS 3.31f
C1707 a_1500_55738# VSUBS 0.625f
C1708 a_n1558_55738# VSUBS 0.625f
C1709 a_n1500_55641# VSUBS 3.31f
C1710 a_1500_56974# VSUBS 0.625f
C1711 a_n1558_56974# VSUBS 0.625f
C1712 a_n1500_56877# VSUBS 3.31f
C1713 a_1500_58210# VSUBS 0.625f
C1714 a_n1558_58210# VSUBS 0.625f
C1715 a_n1500_58113# VSUBS 3.31f
C1716 a_1500_59446# VSUBS 0.625f
C1717 a_n1558_59446# VSUBS 0.625f
C1718 a_n1500_59349# VSUBS 3.31f
C1719 a_1500_60682# VSUBS 0.625f
C1720 a_n1558_60682# VSUBS 0.625f
C1721 a_n1500_60585# VSUBS 3.31f
C1722 a_1500_61918# VSUBS 0.638f
C1723 a_n1558_61918# VSUBS 0.638f
C1724 a_n1500_61821# VSUBS 5.03f
C1725 w_n1594_n63018# VSUBS 11.5f
C1726 w_n1594_n61782# VSUBS 11.5f
C1727 w_n1594_n60546# VSUBS 11.5f
C1728 w_n1594_n59310# VSUBS 11.5f
C1729 w_n1594_n58074# VSUBS 11.5f
C1730 w_n1594_n56838# VSUBS 11.5f
C1731 w_n1594_n55602# VSUBS 11.5f
C1732 w_n1594_n54366# VSUBS 11.5f
C1733 w_n1594_n53130# VSUBS 11.5f
C1734 w_n1594_n51894# VSUBS 11.5f
C1735 w_n1594_n50658# VSUBS 11.5f
C1736 w_n1594_n49422# VSUBS 11.5f
C1737 w_n1594_n48186# VSUBS 11.5f
C1738 w_n1594_n46950# VSUBS 11.5f
C1739 w_n1594_n45714# VSUBS 11.5f
C1740 w_n1594_n44478# VSUBS 11.5f
C1741 w_n1594_n43242# VSUBS 11.5f
C1742 w_n1594_n42006# VSUBS 11.5f
C1743 w_n1594_n40770# VSUBS 11.5f
C1744 w_n1594_n39534# VSUBS 11.5f
C1745 w_n1594_n38298# VSUBS 11.5f
C1746 w_n1594_n37062# VSUBS 11.5f
C1747 w_n1594_n35826# VSUBS 11.5f
C1748 w_n1594_n34590# VSUBS 11.5f
C1749 w_n1594_n33354# VSUBS 11.5f
C1750 w_n1594_n32118# VSUBS 11.5f
C1751 w_n1594_n30882# VSUBS 11.5f
C1752 w_n1594_n29646# VSUBS 11.5f
C1753 w_n1594_n28410# VSUBS 11.5f
C1754 w_n1594_n27174# VSUBS 11.5f
C1755 w_n1594_n25938# VSUBS 11.5f
C1756 w_n1594_n24702# VSUBS 11.5f
C1757 w_n1594_n23466# VSUBS 11.5f
C1758 w_n1594_n22230# VSUBS 11.5f
C1759 w_n1594_n20994# VSUBS 11.5f
C1760 w_n1594_n19758# VSUBS 11.5f
C1761 w_n1594_n18522# VSUBS 11.5f
C1762 w_n1594_n17286# VSUBS 11.5f
C1763 w_n1594_n16050# VSUBS 11.5f
C1764 w_n1594_n14814# VSUBS 11.5f
C1765 w_n1594_n13578# VSUBS 11.5f
C1766 w_n1594_n12342# VSUBS 11.5f
C1767 w_n1594_n11106# VSUBS 11.5f
C1768 w_n1594_n9870# VSUBS 11.5f
C1769 w_n1594_n8634# VSUBS 11.5f
C1770 w_n1594_n7398# VSUBS 11.5f
C1771 w_n1594_n6162# VSUBS 11.5f
C1772 w_n1594_n4926# VSUBS 11.5f
C1773 w_n1594_n3690# VSUBS 11.5f
C1774 w_n1594_n2454# VSUBS 11.5f
C1775 w_n1594_n1218# VSUBS 11.5f
C1776 w_n1594_18# VSUBS 11.5f
C1777 w_n1594_1254# VSUBS 11.5f
C1778 w_n1594_2490# VSUBS 11.5f
C1779 w_n1594_3726# VSUBS 11.5f
C1780 w_n1594_4962# VSUBS 11.5f
C1781 w_n1594_6198# VSUBS 11.5f
C1782 w_n1594_7434# VSUBS 11.5f
C1783 w_n1594_8670# VSUBS 11.5f
C1784 w_n1594_9906# VSUBS 11.5f
C1785 w_n1594_11142# VSUBS 11.5f
C1786 w_n1594_12378# VSUBS 11.5f
C1787 w_n1594_13614# VSUBS 11.5f
C1788 w_n1594_14850# VSUBS 11.5f
C1789 w_n1594_16086# VSUBS 11.5f
C1790 w_n1594_17322# VSUBS 11.5f
C1791 w_n1594_18558# VSUBS 11.5f
C1792 w_n1594_19794# VSUBS 11.5f
C1793 w_n1594_21030# VSUBS 11.5f
C1794 w_n1594_22266# VSUBS 11.5f
C1795 w_n1594_23502# VSUBS 11.5f
C1796 w_n1594_24738# VSUBS 11.5f
C1797 w_n1594_25974# VSUBS 11.5f
C1798 w_n1594_27210# VSUBS 11.5f
C1799 w_n1594_28446# VSUBS 11.5f
C1800 w_n1594_29682# VSUBS 11.5f
C1801 w_n1594_30918# VSUBS 11.5f
C1802 w_n1594_32154# VSUBS 11.5f
C1803 w_n1594_33390# VSUBS 11.5f
C1804 w_n1594_34626# VSUBS 11.5f
C1805 w_n1594_35862# VSUBS 11.5f
C1806 w_n1594_37098# VSUBS 11.5f
C1807 w_n1594_38334# VSUBS 11.5f
C1808 w_n1594_39570# VSUBS 11.5f
C1809 w_n1594_40806# VSUBS 11.5f
C1810 w_n1594_42042# VSUBS 11.5f
C1811 w_n1594_43278# VSUBS 11.5f
C1812 w_n1594_44514# VSUBS 11.5f
C1813 w_n1594_45750# VSUBS 11.5f
C1814 w_n1594_46986# VSUBS 11.5f
C1815 w_n1594_48222# VSUBS 11.5f
C1816 w_n1594_49458# VSUBS 11.5f
C1817 w_n1594_50694# VSUBS 11.5f
C1818 w_n1594_51930# VSUBS 11.5f
C1819 w_n1594_53166# VSUBS 11.5f
C1820 w_n1594_54402# VSUBS 11.5f
C1821 w_n1594_55638# VSUBS 11.5f
C1822 w_n1594_56874# VSUBS 11.5f
C1823 w_n1594_58110# VSUBS 11.5f
C1824 w_n1594_59346# VSUBS 11.5f
C1825 w_n1594_60582# VSUBS 11.5f
C1826 w_n1594_61818# VSUBS 11.5f
.ends

.subckt sky130_fd_pr__pfet_01v8_UDMRD5 a_n558_n10388# a_n558_n7916# a_n500_5583# a_n500_n10485#
+ a_500_1972# a_n558_8152# a_n500_8055# a_500_4444# w_n594_3108# w_n594_6816# a_500_n2972#
+ a_500_736# a_500_n5444# a_n500_n597# w_n594_636# a_500_n500# a_500_9388# w_n594_n3072#
+ a_n558_1972# w_n594_n6780# w_n594_n600# a_n500_1875# a_n558_4444# w_n594_n9252#
+ a_n500_4347# a_n558_n6680# w_n594_n10488# a_n558_n9152# a_n500_n5541# a_n500_639#
+ a_500_3208# a_n500_n8013# a_500_6916# a_500_n1736# a_n558_n500# a_n558_9388# a_500_n4208#
+ w_n594_5580# a_500_n7916# w_n594_8052# w_n594_n5544# a_n558_736# a_n558_3208# w_n594_n8016#
+ a_n558_n2972# a_n558_6916# a_n558_n5444# a_n500_n1833# a_n500_6819# a_n500_n4305#
+ w_n594_1872# a_500_5680# a_n500_9291# a_n500_n3069# w_n594_4344# a_n500_n6777# a_500_8152#
+ w_n594_n1836# a_n500_n9249# a_500_n6680# w_n594_n4308# a_500_n10388# a_n500_3111#
+ a_500_n9152# a_n558_n1736# w_n594_9288# a_n558_n4208# a_n558_5680# VSUBS
X0 a_500_1972# a_n500_1875# a_n558_1972# w_n594_1872# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X1 a_500_6916# a_n500_6819# a_n558_6916# w_n594_6816# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X2 a_500_4444# a_n500_4347# a_n558_4444# w_n594_4344# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X3 a_500_n9152# a_n500_n9249# a_n558_n9152# w_n594_n9252# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X4 a_500_3208# a_n500_3111# a_n558_3208# w_n594_3108# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X5 a_500_n2972# a_n500_n3069# a_n558_n2972# w_n594_n3072# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X6 a_500_n7916# a_n500_n8013# a_n558_n7916# w_n594_n8016# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X7 a_500_9388# a_n500_9291# a_n558_9388# w_n594_9288# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X8 a_500_n5444# a_n500_n5541# a_n558_n5444# w_n594_n5544# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X9 a_500_n500# a_n500_n597# a_n558_n500# w_n594_n600# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X10 a_500_n1736# a_n500_n1833# a_n558_n1736# w_n594_n1836# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X11 a_500_n4208# a_n500_n4305# a_n558_n4208# w_n594_n4308# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X12 a_500_n10388# a_n500_n10485# a_n558_n10388# w_n594_n10488# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X13 a_500_736# a_n500_639# a_n558_736# w_n594_636# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X14 a_500_n6680# a_n500_n6777# a_n558_n6680# w_n594_n6780# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X15 a_500_5680# a_n500_5583# a_n558_5680# w_n594_5580# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
X16 a_500_8152# a_n500_8055# a_n558_8152# w_n594_8052# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=5
**devattr s=58000,2116 d=58000,2116
C0 a_500_6916# w_n594_8052# 0.0023f
C1 w_n594_n1836# a_n500_n3069# 0.00575f
C2 a_n558_n2972# a_n500_n3069# 0.204f
C3 a_n558_n7916# a_500_n7916# 0.0663f
C4 w_n594_n600# a_n558_n1736# 0.0023f
C5 a_n558_n5444# w_n594_n5544# 0.0187f
C6 w_n594_n6780# a_500_n6680# 0.0187f
C7 w_n594_n3072# a_n558_n1736# 0.0023f
C8 a_500_n500# a_n558_n500# 0.0663f
C9 a_n500_n1833# w_n594_n1836# 0.593f
C10 a_n500_n1833# a_n500_n597# 1.03f
C11 a_n500_n4305# w_n594_n4308# 0.593f
C12 a_500_8152# w_n594_6816# 0.0023f
C13 a_500_n1736# a_n558_n1736# 0.0663f
C14 a_n558_1972# w_n594_1872# 0.0187f
C15 a_n500_3111# w_n594_3108# 0.593f
C16 w_n594_n6780# a_n558_n5444# 0.0023f
C17 w_n594_n1836# a_500_n500# 0.0023f
C18 a_n500_n597# a_500_n500# 0.204f
C19 a_500_9388# w_n594_8052# 0.0023f
C20 a_500_736# a_500_1972# 0.0105f
C21 a_n500_n10485# a_n500_n9249# 1.03f
C22 a_n558_4444# a_n558_5680# 0.0105f
C23 a_n500_8055# w_n594_6816# 0.00575f
C24 a_500_3208# w_n594_1872# 0.0023f
C25 a_500_8152# a_n500_8055# 0.204f
C26 w_n594_n9252# a_n558_n9152# 0.0187f
C27 a_n558_1972# a_n500_1875# 0.204f
C28 w_n594_n10488# a_n500_n9249# 0.00575f
C29 a_500_3208# w_n594_4344# 0.0023f
C30 w_n594_636# a_n558_n500# 0.0023f
C31 a_n500_n5541# w_n594_n5544# 0.593f
C32 w_n594_8052# a_n558_8152# 0.0187f
C33 a_500_5680# a_n558_5680# 0.0663f
C34 w_n594_n6780# a_n500_n8013# 0.00575f
C35 a_500_n9152# w_n594_n10488# 0.0023f
C36 a_n558_736# w_n594_1872# 0.0023f
C37 a_500_736# w_n594_n600# 0.0023f
C38 w_n594_636# a_n500_n597# 0.00575f
C39 a_n500_n5541# w_n594_n6780# 0.00575f
C40 w_n594_n8016# a_n558_n6680# 0.0023f
C41 a_n558_n4208# w_n594_n5544# 0.0023f
C42 w_n594_636# a_n500_639# 0.593f
C43 a_n558_3208# a_n558_1972# 0.0105f
C44 w_n594_8052# a_n558_6916# 0.0023f
C45 a_500_n4208# a_500_n5444# 0.0105f
C46 a_n500_4347# a_n500_5583# 1.03f
C47 a_500_n10388# w_n594_n9252# 0.0023f
C48 w_n594_n8016# a_n558_n7916# 0.0187f
C49 a_n558_5680# w_n594_6816# 0.0023f
C50 a_n500_n4305# a_n500_n3069# 1.03f
C51 w_n594_n1836# a_n558_n500# 0.0023f
C52 a_n500_n597# a_n558_n500# 0.204f
C53 a_n500_n10485# a_n558_n10388# 0.204f
C54 a_n558_3208# a_500_3208# 0.0663f
C55 a_n500_5583# w_n594_5580# 0.593f
C56 a_n500_9291# a_500_9388# 0.204f
C57 a_n500_n5541# a_n558_n5444# 0.204f
C58 a_n558_4444# w_n594_4344# 0.0187f
C59 w_n594_n3072# a_500_n4208# 0.0023f
C60 w_n594_n8016# a_n500_n6777# 0.00575f
C61 a_n500_n597# w_n594_n1836# 0.00575f
C62 w_n594_n1836# a_n558_n2972# 0.0023f
C63 a_n500_6819# w_n594_8052# 0.00575f
C64 a_n500_9291# w_n594_9288# 0.593f
C65 w_n594_n10488# a_n558_n10388# 0.0187f
C66 a_500_n2972# a_500_n4208# 0.0105f
C67 a_n500_n597# a_n500_639# 1.03f
C68 a_n558_n5444# a_n558_n4208# 0.0105f
C69 a_500_5680# w_n594_4344# 0.0023f
C70 w_n594_n4308# a_500_n5444# 0.0023f
C71 a_n558_n9152# a_n500_n9249# 0.204f
C72 a_n500_n4305# w_n594_n5544# 0.00575f
C73 a_500_6916# w_n594_5580# 0.0023f
C74 a_n500_n1833# a_n558_n1736# 0.204f
C75 w_n594_n9252# a_n500_n8013# 0.00575f
C76 w_n594_n3072# a_500_n2972# 0.0187f
C77 a_n500_4347# w_n594_5580# 0.00575f
C78 w_n594_n600# a_500_n1736# 0.0023f
C79 a_500_n9152# a_n558_n9152# 0.0663f
C80 w_n594_n4308# a_500_n4208# 0.0187f
C81 a_500_n7916# w_n594_n6780# 0.0023f
C82 a_n558_1972# a_500_1972# 0.0663f
C83 w_n594_n3072# a_500_n1736# 0.0023f
C84 a_500_4444# w_n594_4344# 0.0187f
C85 a_n500_1875# w_n594_3108# 0.00575f
C86 a_500_n2972# a_500_n1736# 0.0105f
C87 a_500_n7916# a_500_n6680# 0.0105f
C88 a_n558_n2972# a_n558_n4208# 0.0105f
C89 a_n558_4444# a_n558_3208# 0.0105f
C90 a_500_n2972# w_n594_n4308# 0.0023f
C91 a_500_3208# a_500_1972# 0.0105f
C92 a_n558_736# a_500_736# 0.0663f
C93 a_n558_n7916# a_n558_n6680# 0.0105f
C94 a_n558_3208# w_n594_3108# 0.0187f
C95 a_500_n9152# a_500_n10388# 0.0105f
C96 w_n594_636# a_n500_1875# 0.00575f
C97 a_500_8152# w_n594_8052# 0.0187f
C98 a_n500_3111# w_n594_1872# 0.00575f
C99 a_n500_3111# w_n594_4344# 0.00575f
C100 a_500_9388# w_n594_9288# 0.0187f
C101 a_n500_n6777# a_n558_n6680# 0.204f
C102 a_n558_n9152# a_n558_n10388# 0.0105f
C103 a_n500_5583# a_n500_6819# 1.03f
C104 a_500_6916# a_n558_6916# 0.0663f
C105 w_n594_n8016# a_n558_n9152# 0.0023f
C106 a_500_n7916# a_n500_n8013# 0.204f
C107 a_n500_639# w_n594_1872# 0.00575f
C108 a_n500_3111# a_n500_1875# 1.03f
C109 a_n500_8055# w_n594_8052# 0.593f
C110 a_500_736# a_500_n500# 0.0105f
C111 a_n558_736# w_n594_n600# 0.0023f
C112 a_n558_n1736# a_n558_n500# 0.0105f
C113 a_n500_n8013# a_n500_n9249# 1.03f
C114 w_n594_n9252# a_500_n7916# 0.0023f
C115 w_n594_5580# a_n558_6916# 0.0023f
C116 w_n594_9288# a_n558_8152# 0.0023f
C117 a_n558_5680# w_n594_4344# 0.0023f
C118 a_n500_n5541# a_n500_n4305# 1.03f
C119 a_n500_1875# a_n500_639# 1.03f
C120 a_500_6916# a_n500_6819# 0.204f
C121 w_n594_n1836# a_n558_n1736# 0.0187f
C122 a_500_n10388# a_n558_n10388# 0.0663f
C123 a_n500_5583# a_500_5680# 0.204f
C124 w_n594_n10488# a_n500_n10485# 0.593f
C125 a_n558_n2972# a_n558_n1736# 0.0105f
C126 w_n594_n9252# a_n500_n9249# 0.593f
C127 a_n558_3208# a_n500_3111# 0.204f
C128 w_n594_n8016# a_500_n6680# 0.0023f
C129 a_500_1972# w_n594_3108# 0.0023f
C130 w_n594_n3072# a_n500_n3069# 0.593f
C131 a_500_n9152# w_n594_n9252# 0.0187f
C132 a_n558_9388# w_n594_8052# 0.0023f
C133 a_500_n2972# a_n500_n3069# 0.204f
C134 a_n500_n1833# w_n594_n600# 0.00575f
C135 a_n500_n4305# a_n558_n4208# 0.204f
C136 w_n594_n5544# a_500_n5444# 0.0187f
C137 a_n500_6819# w_n594_5580# 0.00575f
C138 w_n594_636# a_500_736# 0.0187f
C139 w_n594_n3072# a_n500_n1833# 0.00575f
C140 a_n558_4444# a_n500_4347# 0.204f
C141 a_n558_8152# a_n558_6916# 0.0105f
C142 a_500_n4208# w_n594_n5544# 0.0023f
C143 w_n594_n600# a_500_n500# 0.0187f
C144 a_n500_5583# w_n594_6816# 0.00575f
C145 a_500_6916# a_500_5680# 0.0105f
C146 w_n594_n6780# a_500_n5444# 0.0023f
C147 w_n594_n4308# a_n500_n3069# 0.00575f
C148 a_n500_n1833# a_500_n1736# 0.204f
C149 w_n594_636# a_500_1972# 0.0023f
C150 a_n500_4347# w_n594_3108# 0.00575f
C151 a_n558_4444# w_n594_5580# 0.0023f
C152 a_n558_736# a_n558_1972# 0.0105f
C153 a_500_n6680# a_500_n5444# 0.0105f
C154 a_n500_9291# a_n500_8055# 1.03f
C155 a_500_n500# a_500_n1736# 0.0105f
C156 w_n594_n8016# a_n500_n8013# 0.593f
C157 a_500_5680# w_n594_5580# 0.0187f
C158 a_n500_4347# a_500_4444# 0.204f
C159 a_n558_n6680# w_n594_n5544# 0.0023f
C160 a_n558_n5444# a_500_n5444# 0.0663f
C161 a_500_6916# w_n594_6816# 0.0187f
C162 a_500_8152# a_500_6916# 0.0105f
C163 w_n594_n9252# a_n558_n10388# 0.0023f
C164 a_n558_n7916# a_n558_n9152# 0.0105f
C165 a_500_736# a_n500_639# 0.204f
C166 a_n500_1875# w_n594_1872# 0.593f
C167 a_500_n9152# a_500_n7916# 0.0105f
C168 a_500_4444# w_n594_5580# 0.0023f
C169 w_n594_n6780# a_n558_n6680# 0.0187f
C170 a_n500_9291# a_n558_9388# 0.204f
C171 a_n500_6819# a_n558_6916# 0.204f
C172 a_n558_n6680# a_500_n6680# 0.0663f
C173 a_n558_n7916# w_n594_n6780# 0.0023f
C174 a_500_n9152# a_n500_n9249# 0.204f
C175 a_n500_n6777# w_n594_n5544# 0.00575f
C176 w_n594_n10488# a_n558_n9152# 0.0023f
C177 w_n594_n600# a_n558_n500# 0.0187f
C178 a_n558_1972# w_n594_3108# 0.0023f
C179 a_n558_3208# w_n594_1872# 0.0023f
C180 a_n500_4347# a_n500_3111# 1.03f
C181 a_500_8152# a_500_9388# 0.0105f
C182 a_n500_5583# a_n558_5680# 0.204f
C183 a_n558_n5444# a_n558_n6680# 0.0105f
C184 a_n558_3208# w_n594_4344# 0.0023f
C185 a_n500_n5541# a_500_n5444# 0.204f
C186 a_500_8152# w_n594_9288# 0.0023f
C187 a_n500_n6777# w_n594_n6780# 0.593f
C188 a_n500_n597# w_n594_n600# 0.593f
C189 a_500_n10388# a_n500_n10485# 0.204f
C190 a_n558_n5444# w_n594_n4308# 0.0023f
C191 a_500_3208# w_n594_3108# 0.0187f
C192 w_n594_n600# a_n500_639# 0.00575f
C193 w_n594_n3072# a_n558_n2972# 0.0187f
C194 w_n594_6816# a_n558_8152# 0.0023f
C195 a_n500_n6777# a_500_n6680# 0.204f
C196 a_500_8152# a_n558_8152# 0.0663f
C197 a_500_n2972# w_n594_n1836# 0.0023f
C198 a_500_n2972# a_n558_n2972# 0.0663f
C199 w_n594_636# a_n558_1972# 0.0023f
C200 a_n500_n1833# a_n500_n3069# 1.03f
C201 w_n594_n1836# a_500_n1736# 0.0187f
C202 w_n594_n8016# a_500_n7916# 0.0187f
C203 a_500_n10388# w_n594_n10488# 0.0187f
C204 a_500_4444# a_500_3208# 0.0105f
C205 a_n500_8055# w_n594_9288# 0.00575f
C206 a_500_n4208# a_n558_n4208# 0.0663f
C207 a_500_736# w_n594_1872# 0.0023f
C208 a_n558_n2972# w_n594_n4308# 0.0023f
C209 w_n594_6816# a_n558_6916# 0.0187f
C210 a_n558_n7916# a_n500_n8013# 0.204f
C211 a_n500_8055# a_n558_8152# 0.204f
C212 w_n594_n8016# a_n500_n9249# 0.00575f
C213 a_n558_5680# w_n594_5580# 0.0187f
C214 w_n594_n3072# a_n558_n4208# 0.0023f
C215 w_n594_n8016# a_500_n9152# 0.0023f
C216 a_n558_9388# a_500_9388# 0.0663f
C217 a_500_1972# w_n594_1872# 0.0187f
C218 a_n500_n5541# w_n594_n4308# 0.00575f
C219 w_n594_n9252# a_n558_n7916# 0.0023f
C220 a_n500_5583# w_n594_4344# 0.00575f
C221 w_n594_636# a_n558_736# 0.0187f
C222 a_n500_n6777# a_n500_n8013# 1.03f
C223 a_n558_9388# w_n594_9288# 0.0187f
C224 a_n558_4444# w_n594_3108# 0.0023f
C225 a_500_3208# a_n500_3111# 0.204f
C226 a_n500_6819# w_n594_6816# 0.593f
C227 a_n500_9291# w_n594_8052# 0.00575f
C228 w_n594_n9252# a_n500_n10485# 0.00575f
C229 w_n594_n4308# a_n558_n4208# 0.0187f
C230 a_n558_9388# a_n558_8152# 0.0105f
C231 a_n500_1875# a_500_1972# 0.204f
C232 a_n500_n5541# a_n500_n6777# 1.03f
C233 a_n558_4444# a_500_4444# 0.0663f
C234 a_n558_736# a_n558_n500# 0.0105f
C235 a_n500_n4305# a_500_n4208# 0.204f
C236 a_n500_4347# w_n594_4344# 0.593f
C237 a_500_4444# a_500_5680# 0.0105f
C238 a_n500_8055# a_n500_6819# 1.03f
C239 a_500_4444# w_n594_3108# 0.0023f
C240 w_n594_636# a_500_n500# 0.0023f
C241 a_500_5680# w_n594_6816# 0.0023f
C242 w_n594_n3072# a_n500_n4305# 0.00575f
C243 a_n558_736# a_n500_639# 0.204f
C244 a_500_n6680# w_n594_n5544# 0.0023f
C245 a_n558_5680# a_n558_6916# 0.0105f
C246 a_500_n10388# VSUBS 0.561f
C247 a_n558_n10388# VSUBS 0.561f
C248 a_n500_n10485# VSUBS 1.74f
C249 a_500_n9152# VSUBS 0.548f
C250 a_n558_n9152# VSUBS 0.548f
C251 a_n500_n9249# VSUBS 1.17f
C252 a_500_n7916# VSUBS 0.548f
C253 a_n558_n7916# VSUBS 0.548f
C254 a_n500_n8013# VSUBS 1.17f
C255 a_500_n6680# VSUBS 0.548f
C256 a_n558_n6680# VSUBS 0.548f
C257 a_n500_n6777# VSUBS 1.17f
C258 a_500_n5444# VSUBS 0.548f
C259 a_n558_n5444# VSUBS 0.548f
C260 a_n500_n5541# VSUBS 1.17f
C261 a_500_n4208# VSUBS 0.548f
C262 a_n558_n4208# VSUBS 0.548f
C263 a_n500_n4305# VSUBS 1.17f
C264 a_500_n2972# VSUBS 0.548f
C265 a_n558_n2972# VSUBS 0.548f
C266 a_n500_n3069# VSUBS 1.17f
C267 a_500_n1736# VSUBS 0.548f
C268 a_n558_n1736# VSUBS 0.548f
C269 a_n500_n1833# VSUBS 1.17f
C270 a_500_n500# VSUBS 0.548f
C271 a_n558_n500# VSUBS 0.548f
C272 a_n500_n597# VSUBS 1.17f
C273 a_500_736# VSUBS 0.548f
C274 a_n558_736# VSUBS 0.548f
C275 a_n500_639# VSUBS 1.17f
C276 a_500_1972# VSUBS 0.548f
C277 a_n558_1972# VSUBS 0.548f
C278 a_n500_1875# VSUBS 1.17f
C279 a_500_3208# VSUBS 0.548f
C280 a_n558_3208# VSUBS 0.548f
C281 a_n500_3111# VSUBS 1.17f
C282 a_500_4444# VSUBS 0.548f
C283 a_n558_4444# VSUBS 0.548f
C284 a_n500_4347# VSUBS 1.17f
C285 a_500_5680# VSUBS 0.548f
C286 a_n558_5680# VSUBS 0.548f
C287 a_n500_5583# VSUBS 1.17f
C288 a_500_6916# VSUBS 0.548f
C289 a_n558_6916# VSUBS 0.548f
C290 a_n500_6819# VSUBS 1.17f
C291 a_500_8152# VSUBS 0.548f
C292 a_n558_8152# VSUBS 0.548f
C293 a_n500_8055# VSUBS 1.17f
C294 a_500_9388# VSUBS 0.561f
C295 a_n558_9388# VSUBS 0.561f
C296 a_n500_9291# VSUBS 1.74f
C297 w_n594_n10488# VSUBS 4.28f
C298 w_n594_n9252# VSUBS 4.28f
C299 w_n594_n8016# VSUBS 4.28f
C300 w_n594_n6780# VSUBS 4.28f
C301 w_n594_n5544# VSUBS 4.28f
C302 w_n594_n4308# VSUBS 4.28f
C303 w_n594_n3072# VSUBS 4.28f
C304 w_n594_n1836# VSUBS 4.28f
C305 w_n594_n600# VSUBS 4.28f
C306 w_n594_636# VSUBS 4.28f
C307 w_n594_1872# VSUBS 4.28f
C308 w_n594_3108# VSUBS 4.28f
C309 w_n594_4344# VSUBS 4.28f
C310 w_n594_5580# VSUBS 4.28f
C311 w_n594_6816# VSUBS 4.28f
C312 w_n594_8052# VSUBS 4.28f
C313 w_n594_9288# VSUBS 4.28f
.ends

.subckt sky130_fd_pr__pfet_01v8_RRU5GE a_n300_n1833# w_n394_n1836# a_n358_n1736# a_300_736#
+ w_n394_636# a_n300_n597# a_300_n500# a_n300_639# w_n394_n600# a_300_n1736# a_n358_n500#
+ a_n358_736# VSUBS
X0 a_300_n500# a_n300_n597# a_n358_n500# w_n394_n600# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=3
**devattr s=58000,2116 d=58000,2116
X1 a_300_736# a_n300_639# a_n358_736# w_n394_636# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=3
**devattr s=58000,2116 d=58000,2116
X2 a_300_n1736# a_n300_n1833# a_n358_n1736# w_n394_n1836# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=3
**devattr s=58000,2116 d=58000,2116
C0 a_n300_639# a_300_736# 0.184f
C1 a_300_n500# a_n300_n597# 0.184f
C2 a_300_n500# w_n394_n1836# 0.0023f
C3 a_n358_n500# w_n394_n600# 0.0187f
C4 w_n394_636# a_n358_736# 0.0187f
C5 a_n358_n500# a_n358_736# 0.0105f
C6 a_n358_n500# a_n358_n1736# 0.0105f
C7 w_n394_n600# a_n300_n597# 0.382f
C8 a_n358_n1736# w_n394_n1836# 0.0187f
C9 a_300_n500# w_n394_n600# 0.0187f
C10 a_300_n1736# w_n394_n1836# 0.0187f
C11 w_n394_636# a_300_736# 0.0187f
C12 w_n394_636# a_n300_639# 0.382f
C13 a_n300_n1833# a_n300_n597# 0.62f
C14 a_n300_n1833# w_n394_n1836# 0.382f
C15 a_300_n500# a_300_n1736# 0.0105f
C16 a_n300_639# a_n300_n597# 0.62f
C17 a_n358_736# w_n394_n600# 0.0023f
C18 w_n394_n600# a_n358_n1736# 0.0023f
C19 a_300_n500# a_300_736# 0.0105f
C20 w_n394_n600# a_300_n1736# 0.0023f
C21 a_n358_n1736# a_300_n1736# 0.107f
C22 a_n300_n1833# w_n394_n600# 0.00346f
C23 a_n358_n500# w_n394_636# 0.0023f
C24 w_n394_n600# a_300_736# 0.0023f
C25 a_n300_639# w_n394_n600# 0.00346f
C26 a_n300_n1833# a_n358_n1736# 0.184f
C27 a_n358_736# a_300_736# 0.107f
C28 a_n300_639# a_n358_736# 0.184f
C29 w_n394_636# a_n300_n597# 0.00346f
C30 a_n300_n1833# a_300_n1736# 0.184f
C31 a_n358_n500# a_n300_n597# 0.184f
C32 a_n358_n500# w_n394_n1836# 0.0023f
C33 a_300_n500# w_n394_636# 0.0023f
C34 a_n300_n597# w_n394_n1836# 0.00346f
C35 a_300_n500# a_n358_n500# 0.107f
C36 a_300_n1736# VSUBS 0.536f
C37 a_n358_n1736# VSUBS 0.536f
C38 a_n300_n1833# VSUBS 1.08f
C39 a_300_n500# VSUBS 0.524f
C40 a_n358_n500# VSUBS 0.524f
C41 a_n300_n597# VSUBS 0.739f
C42 a_300_736# VSUBS 0.536f
C43 a_n358_736# VSUBS 0.536f
C44 a_n300_639# VSUBS 1.08f
C45 w_n394_n1836# VSUBS 2.84f
C46 w_n394_n600# VSUBS 2.84f
C47 w_n394_636# VSUBS 2.84f
.ends

.subckt sky130_fd_pr__pfet_01v8_SLZ774 w_n1594_n600# a_n1500_n597# a_1500_n500# a_n1558_n500#
+ VSUBS
X0 a_1500_n500# a_n1500_n597# a_n1558_n500# w_n1594_n600# sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=15
**devattr s=58000,2116 d=58000,2116
C0 w_n1594_n600# a_n1558_n500# 0.0187f
C1 w_n1594_n600# a_1500_n500# 0.0187f
C2 a_n1500_n597# w_n1594_n600# 1.65f
C3 a_n1500_n597# a_n1558_n500# 0.217f
C4 a_n1500_n597# a_1500_n500# 0.217f
C5 a_1500_n500# VSUBS 0.65f
C6 a_n1558_n500# VSUBS 0.65f
C7 a_n1500_n597# VSUBS 6.74f
C8 w_n1594_n600# VSUBS 11.5f
.ends

.subckt opamp_cascode IN_P IN_M VCC VSS OUT VB_A VB_B IB
Xsky130_fd_pr__nfet_01v8_SCE452_3 VSS bias21 bias21 VSS sky130_fd_pr__nfet_01v8_SCE452
XXM9_dummy_15 VCC bias1 dummy_9 dummy_9 VSS sky130_fd_pr__pfet_01v8_ZLZ7XS
XXM5_1 VCC IN_M IN_M bias3 VCC VCC m1_44990_37960# m1_44990_37960# m1_44990_37960#
+ bias3 IN_M bias3 m1_44990_37960# bias3 IN_M m1_44990_37960# bias3 VCC IN_M IN_M
+ bias3 VCC IN_M IN_M IN_M VCC VCC VCC IN_M IN_M IN_M m1_44990_37960# m1_44990_37960#
+ m1_44990_37960# bias3 IN_M VCC bias3 m1_44990_37960# bias3 m1_44990_37960# IN_M
+ VCC bias3 m1_44990_37960# VCC bias3 VCC VCC m1_44990_37960# bias3 m1_44990_37960#
+ bias3 bias3 m1_44990_37960# bias3 VCC m1_44990_37960# IN_M VCC VSS sky130_fd_pr__pfet_01v8_7DHACV
XXM4_dummy_2 dummy_4 bias3 dummy_4 dummy_4 bias3 dummy_4 bias3 dummy_4 bias3 dummy_4
+ dummy_4 dummy_4 dummy_4 dummy_4 bias3 dummy_4 dummy_4 bias3 VSS sky130_fd_pr__nfet_01v8_MHE452
XXM9_dummy_16 VCC bias1 dummy_9 dummy_9 VSS sky130_fd_pr__pfet_01v8_ZLZ7XS
XXM100_4 IB VCC IB IB VCC VCC VCC IB VSS sky130_fd_pr__pfet_01v8_P2UXFR
XXM4_dummy_3 dummy_4 bias3 dummy_4 VSS sky130_fd_pr__nfet_01v8_SCE452
XXM9_dummy_17 VCC bias1 dummy_9 dummy_9 VSS sky130_fd_pr__pfet_01v8_ZLZ7XS
XXM5_dummy_10 dummy_5 IN_P VCC dummy_5 VSS sky130_fd_pr__pfet_01v8_MGA63L
XXM9_dummy_18 VCC bias1 dummy_9 dummy_9 VSS sky130_fd_pr__pfet_01v8_ZLZ7XS
Xsky130_fd_pr__nfet_01v8_VT3ZQW_0 dummy_4 bias3 dummy_4 VSS sky130_fd_pr__nfet_01v8_VT3ZQW
XXM9_dummy_19 VCC bias1 dummy_9 dummy_9 VSS sky130_fd_pr__pfet_01v8_ZLZ7XS
Xsky130_fd_pr__pfet_01v8_RRUZAE_0 dummy_100 IB IB VCC VCC dummy_100 dummy_100 dummy_100
+ dummy_100 VCC VCC IB dummy_100 IB dummy_100 IB VCC dummy_100 dummy_100 dummy_100
+ VSS sky130_fd_pr__pfet_01v8_RRUZAE
Xsky130_fd_pr__pfet_01v8_P2UXFR_0 IB VCC VCC IB IB VCC IB VCC VSS sky130_fd_pr__pfet_01v8_P2UXFR
XXM4_dummy_7 dummy_4 bias3 dummy_4 VSS sky130_fd_pr__nfet_01v8_SCE452
Xsky130_fd_pr__pfet_01v8_ZLZ7XS_0 VCC bias1 dummy_9 dummy_9 VSS sky130_fd_pr__pfet_01v8_ZLZ7XS
Xsky130_fd_pr__pfet_01v8_8DHNHY_0 VCC IN_P IN_P dummy_5 IN_P VCC dummy_5 VCC dummy_5
+ dummy_5 dummy_5 dummy_5 IN_P dummy_5 dummy_5 VCC dummy_5 IN_P dummy_5 dummy_5 VCC
+ dummy_5 IN_P IN_P dummy_5 VCC IN_P IN_P IN_P VCC VCC dummy_5 VCC IN_P IN_P VCC IN_P
+ dummy_5 dummy_5 dummy_5 dummy_5 IN_P VCC dummy_5 dummy_5 dummy_5 dummy_5 IN_P VCC
+ dummy_5 dummy_5 VCC dummy_5 dummy_5 VCC VCC dummy_5 dummy_5 dummy_5 dummy_5 dummy_5
+ dummy_5 dummy_5 VCC IN_P dummy_5 IN_P VCC VSS sky130_fd_pr__pfet_01v8_8DHNHY
XXM100_dummy_1 dummy_100 IB IB VCC VCC dummy_100 dummy_100 dummy_100 dummy_100 VCC
+ VCC IB dummy_100 IB dummy_100 IB VCC dummy_100 dummy_100 dummy_100 VSS sky130_fd_pr__pfet_01v8_RRUZAE
XXM1_1 m1m2 m1m2 bias1 VCC bias1 m1m2 VCC bias1 VCC VCC VCC bias1 m1m2 VCC VCC m1m2
+ VCC bias1 bias1 VCC VCC VCC bias1 m1m2 m1m2 m1m2 m1m2 bias1 VCC m1m2 VCC bias1 VCC
+ VCC VCC m1m2 m1m2 VCC bias1 VCC bias1 m1m2 bias1 VCC m1m2 VCC bias1 m1m2 VCC bias1
+ m1m2 VCC VCC VCC VCC VCC bias1 VCC VCC bias1 m1m2 m1m2 bias1 bias1 VCC VCC VCC m1m2
+ bias1 VCC bias1 VCC m1m2 VCC bias1 m1m2 VCC VCC VCC VCC VCC m1m2 VCC m1m2 bias1
+ m1m2 bias1 VCC bias1 bias1 bias1 VCC VCC VCC bias1 m1m2 VCC m1m2 VCC bias1 m1m2
+ m1m2 VCC VCC bias1 VCC m1m2 m1m2 VCC bias1 VCC m1m2 m1m2 bias1 VCC bias1 VCC VCC
+ m1m2 m1m2 VCC bias1 VCC VCC m1m2 VCC bias1 bias1 VCC VCC m1m2 VCC bias1 m1m2 VCC
+ m1m2 bias1 VCC VCC VCC m1m2 m1m2 VCC VCC VCC VCC VCC bias1 bias1 m1m2 m1m2 VCC m1m2
+ VCC VCC m1m2 VCC VCC VCC bias1 VCC m1m2 bias1 VCC VCC m1m2 m1m2 m1m2 VCC VCC m1m2
+ VCC VCC VCC m1m2 bias1 m1m2 bias1 bias1 VCC bias1 VCC VCC bias1 VCC bias1 VCC m1m2
+ VCC m1m2 m1m2 bias1 bias1 VCC bias1 bias1 VCC bias1 VCC m1m2 m1m2 VCC bias1 bias1
+ VCC VCC m1m2 m1m2 bias1 VCC bias1 VCC VCC VCC VCC bias1 m1m2 m1m2 bias1 m1m2 bias1
+ VCC VCC VCC VCC bias1 m1m2 m1m2 VCC bias1 bias1 VCC VCC bias1 VCC VCC m1m2 bias1
+ VCC VCC VCC bias1 m1m2 bias1 VCC bias1 VCC VCC bias1 VCC VCC VCC bias1 VCC bias1
+ m1m2 m1m2 VCC VCC VCC VCC bias1 VCC VCC VCC VCC VCC m1m2 bias1 bias1 VCC m1m2 VCC
+ VCC VCC bias1 bias1 VCC VCC VCC VCC m1m2 m1m2 m1m2 VCC VCC VCC VCC bias1 VCC VCC
+ m1m2 bias1 VCC VCC VCC bias1 bias1 VCC VCC m1m2 m1m2 bias1 m1m2 VCC VCC bias1 m1m2
+ VCC bias1 m1m2 m1m2 VCC VCC m1m2 VCC VCC m1m2 VCC bias1 m1m2 m1m2 bias1 m1m2 VCC
+ bias1 VCC VCC bias1 VCC bias1 VCC VCC bias1 VCC VCC VCC m1m2 VCC VCC VCC bias1 VCC
+ m1m2 VCC bias1 m1m2 VCC m1m2 m1m2 m1m2 VCC bias1 m1m2 VCC VCC VCC VCC bias1 VCC
+ bias1 m1m2 VCC m1m2 VCC m1m2 VCC VCC VCC bias1 VCC bias1 bias1 m1m2 bias1 VCC VCC
+ VCC VCC VCC VCC VCC VCC bias1 VCC VCC m1m2 bias1 VCC VCC bias1 VCC m1m2 m1m2 VCC
+ m1m2 VCC VCC VSS VCC m1m2 sky130_fd_pr__pfet_01v8_F76D73
XXM4_dummy_9 dummy_4 bias3 dummy_4 VSS sky130_fd_pr__nfet_01v8_SCE452
XXM1_2 m1m2 m1m2 bias1 VCC bias1 m1m2 VCC bias1 VCC VCC VCC bias1 m1m2 VCC VCC m1m2
+ VCC bias1 bias1 VCC VCC VCC bias1 m1m2 m1m2 m1m2 m1m2 bias1 VCC m1m2 VCC bias1 VCC
+ VCC VCC m1m2 m1m2 VCC bias1 VCC bias1 m1m2 bias1 VCC m1m2 VCC bias1 m1m2 VCC bias1
+ m1m2 VCC VCC VCC VCC VCC bias1 VCC VCC bias1 m1m2 m1m2 bias1 bias1 VCC VCC VCC m1m2
+ bias1 VCC bias1 VCC m1m2 VCC bias1 m1m2 VCC VCC VCC VCC VCC m1m2 VCC m1m2 bias1
+ m1m2 bias1 VCC bias1 bias1 bias1 VCC VCC VCC bias1 m1m2 VCC m1m2 VCC bias1 m1m2
+ m1m2 VCC VCC bias1 VCC m1m2 m1m2 VCC bias1 VCC m1m2 m1m2 bias1 VCC bias1 VCC VCC
+ m1m2 m1m2 VCC bias1 VCC VCC m1m2 VCC bias1 bias1 VCC VCC m1m2 VCC bias1 m1m2 VCC
+ m1m2 bias1 VCC VCC VCC m1m2 m1m2 VCC VCC VCC VCC VCC bias1 bias1 m1m2 m1m2 VCC m1m2
+ VCC VCC m1m2 VCC VCC VCC bias1 VCC m1m2 bias1 VCC VCC m1m2 m1m2 m1m2 VCC VCC m1m2
+ VCC VCC VCC m1m2 bias1 m1m2 bias1 bias1 VCC bias1 VCC VCC bias1 VCC bias1 VCC m1m2
+ VCC m1m2 m1m2 bias1 bias1 VCC bias1 bias1 VCC bias1 VCC m1m2 m1m2 VCC bias1 bias1
+ VCC VCC m1m2 m1m2 bias1 VCC bias1 VCC VCC VCC VCC bias1 m1m2 m1m2 bias1 m1m2 bias1
+ VCC VCC VCC VCC bias1 m1m2 m1m2 VCC bias1 bias1 VCC VCC bias1 VCC VCC m1m2 bias1
+ VCC VCC VCC bias1 m1m2 bias1 VCC bias1 VCC VCC bias1 VCC VCC VCC bias1 VCC bias1
+ m1m2 m1m2 VCC VCC VCC VCC bias1 VCC VCC VCC VCC VCC m1m2 bias1 bias1 VCC m1m2 VCC
+ VCC VCC bias1 bias1 VCC VCC VCC VCC m1m2 m1m2 m1m2 VCC VCC VCC VCC bias1 VCC VCC
+ m1m2 bias1 VCC VCC VCC bias1 bias1 VCC VCC m1m2 m1m2 bias1 m1m2 VCC VCC bias1 m1m2
+ VCC bias1 m1m2 m1m2 VCC VCC m1m2 VCC VCC m1m2 VCC bias1 m1m2 m1m2 bias1 m1m2 VCC
+ bias1 VCC VCC bias1 VCC bias1 VCC VCC bias1 VCC VCC VCC m1m2 VCC VCC VCC bias1 VCC
+ m1m2 VCC bias1 m1m2 VCC m1m2 m1m2 m1m2 VCC bias1 m1m2 VCC VCC VCC VCC bias1 VCC
+ bias1 m1m2 VCC m1m2 VCC m1m2 VCC VCC VCC bias1 VCC bias1 bias1 m1m2 bias1 VCC VCC
+ VCC VCC VCC VCC VCC VCC bias1 VCC VCC m1m2 bias1 VCC VCC bias1 VCC m1m2 m1m2 VCC
+ m1m2 VCC VCC VSS VCC m1m2 sky130_fd_pr__pfet_01v8_F76D73
XXM3_dummy_1 VB_B dummy_3 dummy_3 dummy_3 VB_B dummy_3 VB_B VB_B VB_B VB_B dummy_3
+ dummy_3 dummy_3 dummy_3 dummy_3 dummy_3 VB_B dummy_3 dummy_3 dummy_3 VB_B dummy_3
+ dummy_3 dummy_3 VB_B dummy_3 dummy_3 dummy_3 dummy_3 VB_B dummy_3 dummy_3 VB_B VB_B
+ dummy_3 dummy_3 VB_B dummy_3 VB_B dummy_3 VB_B VB_B dummy_3 VB_B dummy_3 dummy_3
+ dummy_3 dummy_3 dummy_3 dummy_3 dummy_3 VSS sky130_fd_pr__nfet_01v8_WK8VRD
XXM100_dummy_3 IB VCC dummy_100 IB dummy_100 VCC dummy_100 dummy_100 VSS sky130_fd_pr__pfet_01v8_P2UXFR
XXM1_3 m1m2 m1m2 bias1 VCC bias1 m1m2 VCC bias1 VCC VCC VCC bias1 m1m2 VCC VCC m1m2
+ VCC bias1 bias1 VCC VCC VCC bias1 m1m2 m1m2 m1m2 m1m2 bias1 VCC m1m2 VCC bias1 VCC
+ VCC VCC m1m2 m1m2 VCC bias1 VCC bias1 m1m2 bias1 VCC m1m2 VCC bias1 m1m2 VCC bias1
+ m1m2 VCC VCC VCC VCC VCC bias1 VCC VCC bias1 m1m2 m1m2 bias1 bias1 VCC VCC VCC m1m2
+ bias1 VCC bias1 VCC m1m2 VCC bias1 m1m2 VCC VCC VCC VCC VCC m1m2 VCC m1m2 bias1
+ m1m2 bias1 VCC bias1 bias1 bias1 VCC VCC VCC bias1 m1m2 VCC m1m2 VCC bias1 m1m2
+ m1m2 VCC VCC bias1 VCC m1m2 m1m2 VCC bias1 VCC m1m2 m1m2 bias1 VCC bias1 VCC VCC
+ m1m2 m1m2 VCC bias1 VCC VCC m1m2 VCC bias1 bias1 VCC VCC m1m2 VCC bias1 m1m2 VCC
+ m1m2 bias1 VCC VCC VCC m1m2 m1m2 VCC VCC VCC VCC VCC bias1 bias1 m1m2 m1m2 VCC m1m2
+ VCC VCC m1m2 VCC VCC VCC bias1 VCC m1m2 bias1 VCC VCC m1m2 m1m2 m1m2 VCC VCC m1m2
+ VCC VCC VCC m1m2 bias1 m1m2 bias1 bias1 VCC bias1 VCC VCC bias1 VCC bias1 VCC m1m2
+ VCC m1m2 m1m2 bias1 bias1 VCC bias1 bias1 VCC bias1 VCC m1m2 m1m2 VCC bias1 bias1
+ VCC VCC m1m2 m1m2 bias1 VCC bias1 VCC VCC VCC VCC bias1 m1m2 m1m2 bias1 m1m2 bias1
+ VCC VCC VCC VCC bias1 m1m2 m1m2 VCC bias1 bias1 VCC VCC bias1 VCC VCC m1m2 bias1
+ VCC VCC VCC bias1 m1m2 bias1 VCC bias1 VCC VCC bias1 VCC VCC VCC bias1 VCC bias1
+ m1m2 m1m2 VCC VCC VCC VCC bias1 VCC VCC VCC VCC VCC m1m2 bias1 bias1 VCC m1m2 VCC
+ VCC VCC bias1 bias1 VCC VCC VCC VCC m1m2 m1m2 m1m2 VCC VCC VCC VCC bias1 VCC VCC
+ m1m2 bias1 VCC VCC VCC bias1 bias1 VCC VCC m1m2 m1m2 bias1 m1m2 VCC VCC bias1 m1m2
+ VCC bias1 m1m2 m1m2 VCC VCC m1m2 VCC VCC m1m2 VCC bias1 m1m2 m1m2 bias1 m1m2 VCC
+ bias1 VCC VCC bias1 VCC bias1 VCC VCC bias1 VCC VCC VCC m1m2 VCC VCC VCC bias1 VCC
+ m1m2 VCC bias1 m1m2 VCC m1m2 m1m2 m1m2 VCC bias1 m1m2 VCC VCC VCC VCC bias1 VCC
+ bias1 m1m2 VCC m1m2 VCC m1m2 VCC VCC VCC bias1 VCC bias1 bias1 m1m2 bias1 VCC VCC
+ VCC VCC VCC VCC VCC VCC bias1 VCC VCC m1m2 bias1 VCC VCC bias1 VCC m1m2 m1m2 VCC
+ m1m2 VCC VCC VSS VCC m1m2 sky130_fd_pr__pfet_01v8_F76D73
XXM100_dummy_4 IB VCC dummy_100 IB dummy_100 VCC dummy_100 dummy_100 VSS sky130_fd_pr__pfet_01v8_P2UXFR
Xsky130_fd_pr__pfet_01v8_MGA63L_0 dummy_5 IN_P VCC dummy_5 VSS sky130_fd_pr__pfet_01v8_MGA63L
XXM3_dummy_3 dummy_3 dummy_3 VB_B VSS sky130_fd_pr__nfet_01v8_AH5E2K
XXM100_dummy_5 IB dummy_100 VCC dummy_100 VSS sky130_fd_pr__pfet_01v8_C2U9V5
XXM1 m1m2 m1m2 bias1 VCC bias1 m1m2 VCC bias1 VCC VCC VCC bias1 m1m2 VCC VCC m1m2
+ VCC bias1 bias1 VCC VCC VCC bias1 m1m2 m1m2 m1m2 m1m2 bias1 VCC m1m2 VCC bias1 VCC
+ VCC VCC m1m2 m1m2 VCC bias1 VCC bias1 m1m2 bias1 VCC m1m2 VCC bias1 m1m2 VCC bias1
+ m1m2 VCC VCC VCC VCC VCC bias1 VCC VCC bias1 m1m2 m1m2 bias1 bias1 VCC VCC VCC m1m2
+ bias1 VCC bias1 VCC m1m2 VCC bias1 m1m2 VCC VCC VCC VCC VCC m1m2 VCC m1m2 bias1
+ m1m2 bias1 VCC bias1 bias1 bias1 VCC VCC VCC bias1 m1m2 VCC m1m2 VCC bias1 m1m2
+ m1m2 VCC VCC bias1 VCC m1m2 m1m2 VCC bias1 VCC m1m2 m1m2 bias1 VCC bias1 VCC VCC
+ m1m2 m1m2 VCC bias1 VCC VCC m1m2 VCC bias1 bias1 VCC VCC m1m2 VCC bias1 m1m2 VCC
+ m1m2 bias1 VCC VCC VCC m1m2 m1m2 VCC VCC VCC VCC VCC bias1 bias1 m1m2 m1m2 VCC m1m2
+ VCC VCC m1m2 VCC VCC VCC bias1 VCC m1m2 bias1 VCC VCC m1m2 m1m2 m1m2 VCC VCC m1m2
+ VCC VCC VCC m1m2 bias1 m1m2 bias1 bias1 VCC bias1 VCC VCC bias1 VCC bias1 VCC m1m2
+ VCC m1m2 m1m2 bias1 bias1 VCC bias1 bias1 VCC bias1 VCC m1m2 m1m2 VCC bias1 bias1
+ VCC VCC m1m2 m1m2 bias1 VCC bias1 VCC VCC VCC VCC bias1 m1m2 m1m2 bias1 m1m2 bias1
+ VCC VCC VCC VCC bias1 m1m2 m1m2 VCC bias1 bias1 VCC VCC bias1 VCC VCC m1m2 bias1
+ VCC VCC VCC bias1 m1m2 bias1 VCC bias1 VCC VCC bias1 VCC VCC VCC bias1 VCC bias1
+ m1m2 m1m2 VCC VCC VCC VCC bias1 VCC VCC VCC VCC VCC m1m2 bias1 bias1 VCC m1m2 VCC
+ VCC VCC bias1 bias1 VCC VCC VCC VCC m1m2 m1m2 m1m2 VCC VCC VCC VCC bias1 VCC VCC
+ m1m2 bias1 VCC VCC VCC bias1 bias1 VCC VCC m1m2 m1m2 bias1 m1m2 VCC VCC bias1 m1m2
+ VCC bias1 m1m2 m1m2 VCC VCC m1m2 VCC VCC m1m2 VCC bias1 m1m2 m1m2 bias1 m1m2 VCC
+ bias1 VCC VCC bias1 VCC bias1 VCC VCC bias1 VCC VCC VCC m1m2 VCC VCC VCC bias1 VCC
+ m1m2 VCC bias1 m1m2 VCC m1m2 m1m2 m1m2 VCC bias1 m1m2 VCC VCC VCC VCC bias1 VCC
+ bias1 m1m2 VCC m1m2 VCC m1m2 VCC VCC VCC bias1 VCC bias1 bias1 m1m2 bias1 VCC VCC
+ VCC VCC VCC VCC VCC VCC bias1 VCC VCC m1m2 bias1 VCC VCC bias1 VCC m1m2 m1m2 VCC
+ m1m2 VCC VCC VSS VCC m1m2 sky130_fd_pr__pfet_01v8_F76D73
XXM100_dummy_6 IB dummy_100 VCC dummy_100 VSS sky130_fd_pr__pfet_01v8_C2U9V5
XXM3_dummy_4 dummy_3 dummy_3 VB_B VSS sky130_fd_pr__nfet_01v8_AH5E2K
Xsky130_fd_pr__nfet_01v8_QP5WRD_0 bias1 bias1 VB_B bias1 VB_B VB_B VB_B VB_B m3m4
+ m3m4 m3m4 m3m4 bias1 bias1 VB_B bias1 bias1 VB_B bias1 bias1 m3m4 VB_B m3m4 m3m4
+ m3m4 m3m4 m3m4 VB_B VB_B bias1 bias1 VB_B bias1 VB_B bias1 VB_B VB_B m3m4 VB_B m3m4
+ m3m4 m3m4 m3m4 bias1 bias1 VSS sky130_fd_pr__nfet_01v8_QP5WRD
XXM2 bias1 VB_A m1m2 bias1 VB_A m1m2 VCC VCC m1m2 m1m2 m1m2 VB_A VCC m1m2 VCC bias1
+ VCC VCC VB_A bias1 VCC VB_A bias1 bias1 VB_A VB_A m1m2 VB_A m1m2 m1m2 bias1 m1m2
+ VCC m1m2 VCC VCC bias1 bias1 VCC bias1 bias1 bias1 VB_A VB_A VB_A VCC m1m2 VB_A
+ VCC VB_A m1m2 VCC VB_A m1m2 VCC VB_A m1m2 bias1 bias1 bias1 VSS sky130_fd_pr__pfet_01v8_UDM5A5
XXM100_dummy_7 IB dummy_100 VCC dummy_100 VSS sky130_fd_pr__pfet_01v8_C2U9V5
XXM4_dummy_10 dummy_4 bias3 dummy_4 VSS sky130_fd_pr__nfet_01v8_SCE452
XXM3 m3m4 m3m4 VB_B m3m4 VB_B VB_B VB_B VB_B bias1 bias1 bias1 bias1 m3m4 m3m4 VB_B
+ m3m4 m3m4 VB_B m3m4 m3m4 bias1 VB_B bias1 bias1 bias1 bias1 bias1 VB_B VB_B m3m4
+ m3m4 VB_B m3m4 VB_B m3m4 VB_B VB_B bias1 VB_B bias1 bias1 bias1 bias1 m3m4 m3m4
+ VSS sky130_fd_pr__nfet_01v8_QP5WRD
XXM8_1 VSS bias21 bias21 VSS sky130_fd_pr__nfet_01v8_VT3ZQW
XXM3_dummy_6 dummy_3 dummy_3 VB_B VSS sky130_fd_pr__nfet_01v8_AH5E2K
XXM100_dummy_8 IB dummy_100 VCC dummy_100 VSS sky130_fd_pr__pfet_01v8_C2U9V5
XXM4 VSS m3m4 bias3 VSS sky130_fd_pr__nfet_01v8_3ZAA45
XXM100_dummy_9 IB dummy_100 VCC dummy_100 VSS sky130_fd_pr__pfet_01v8_C2U9V5
XXM3_dummy_7 dummy_3 dummy_3 VB_B VSS sky130_fd_pr__nfet_01v8_AH5E2K
XXM5 VCC IN_M IN_M m1_44990_37960# VCC VCC bias3 bias3 bias3 m1_44990_37960# IN_M
+ m1_44990_37960# bias3 m1_44990_37960# IN_M bias3 m1_44990_37960# VCC IN_M IN_M m1_44990_37960#
+ VCC IN_M IN_M IN_M VCC VCC VCC IN_M IN_M IN_M bias3 bias3 bias3 m1_44990_37960#
+ IN_M VCC m1_44990_37960# bias3 m1_44990_37960# bias3 IN_M VCC m1_44990_37960# bias3
+ VCC m1_44990_37960# VCC VCC bias3 m1_44990_37960# bias3 m1_44990_37960# m1_44990_37960#
+ bias3 m1_44990_37960# VCC bias3 IN_M VCC VSS sky130_fd_pr__pfet_01v8_7DHACV
XXM8_3 VSS bias21 bias21 VSS sky130_fd_pr__nfet_01v8_VT3ZQW
XXM3_dummy_8 dummy_3 dummy_3 VB_B VSS sky130_fd_pr__nfet_01v8_AH5E2K
XXM6 bias3 bias3 VSS VSS sky130_fd_pr__nfet_01v8_VT3ZQW
XXM3_dummy_9 dummy_3 dummy_3 VB_B VSS sky130_fd_pr__nfet_01v8_AH5E2K
Xsky130_fd_pr__pfet_01v8_SKU9VM_0 VB_A dummy_2 VCC dummy_2 VSS sky130_fd_pr__pfet_01v8_SKU9VM
XXM6_1 bias3 bias3 VSS VSS sky130_fd_pr__nfet_01v8_VT3ZQW
XXM7 VCC IN_P IN_P bias21 VCC VCC m1_44990_37960# m1_44990_37960# m1_44990_37960#
+ bias21 IN_P bias21 m1_44990_37960# bias21 IN_P m1_44990_37960# bias21 VCC IN_P IN_P
+ bias21 VCC IN_P IN_P IN_P VCC VCC VCC IN_P IN_P IN_P m1_44990_37960# m1_44990_37960#
+ m1_44990_37960# bias21 IN_P VCC bias21 m1_44990_37960# bias21 m1_44990_37960# IN_P
+ VCC bias21 m1_44990_37960# VCC bias21 VCC VCC m1_44990_37960# bias21 m1_44990_37960#
+ bias21 bias21 m1_44990_37960# bias21 VCC m1_44990_37960# IN_P VCC VSS sky130_fd_pr__pfet_01v8_7DHACV
Xsky130_fd_pr__pfet_01v8_E769TZ_0 dummy_9 dummy_9 bias1 VCC bias1 dummy_9 dummy_9
+ bias1 VCC VCC dummy_9 bias1 dummy_9 VCC VCC dummy_9 dummy_9 dummy_9 bias1 bias1
+ VCC VCC dummy_9 bias1 dummy_9 dummy_9 dummy_9 dummy_9 bias1 VCC dummy_9 dummy_9
+ bias1 VCC dummy_9 dummy_9 dummy_9 dummy_9 VCC bias1 VCC bias1 dummy_9 bias1 dummy_9
+ dummy_9 dummy_9 bias1 dummy_9 dummy_9 bias1 dummy_9 bias1 VCC VCC dummy_9 VCC VCC
+ bias1 dummy_9 dummy_9 bias1 dummy_9 dummy_9 bias1 bias1 VCC VCC dummy_9 dummy_9
+ bias1 dummy_9 bias1 dummy_9 dummy_9 dummy_9 bias1 dummy_9 VCC VCC dummy_9 VCC VCC
+ dummy_9 VCC dummy_9 bias1 dummy_9 bias1 dummy_9 bias1 bias1 bias1 VCC dummy_9 VCC
+ bias1 dummy_9 dummy_9 dummy_9 dummy_9 bias1 dummy_9 dummy_9 VCC bias1 VCC VCC dummy_9
+ dummy_9 dummy_9 bias1 dummy_9 dummy_9 dummy_9 bias1 VCC bias1 dummy_9 VCC dummy_9
+ dummy_9 dummy_9 VCC bias1 VCC dummy_9 dummy_9 dummy_9 bias1 bias1 dummy_9 dummy_9
+ dummy_9 dummy_9 VCC bias1 dummy_9 VCC dummy_9 bias1 VCC dummy_9 VCC dummy_9 dummy_9
+ dummy_9 VCC VCC dummy_9 VCC VCC bias1 bias1 dummy_9 dummy_9 dummy_9 dummy_9 dummy_9
+ dummy_9 dummy_9 VCC VCC dummy_9 dummy_9 bias1 dummy_9 dummy_9 bias1 VCC dummy_9
+ dummy_9 dummy_9 dummy_9 VCC dummy_9 dummy_9 dummy_9 VCC VCC dummy_9 bias1 dummy_9
+ bias1 bias1 dummy_9 bias1 VCC dummy_9 bias1 VCC bias1 VCC dummy_9 VCC dummy_9 dummy_9
+ bias1 bias1 dummy_9 bias1 bias1 VCC bias1 dummy_9 dummy_9 dummy_9 VCC bias1 bias1
+ VCC VCC dummy_9 dummy_9 bias1 dummy_9 bias1 dummy_9 dummy_9 VCC bias1 dummy_9 bias1
+ dummy_9 dummy_9 bias1 dummy_9 bias1 VCC dummy_9 dummy_9 dummy_9 bias1 dummy_9 dummy_9
+ dummy_9 bias1 bias1 dummy_9 dummy_9 bias1 VCC dummy_9 dummy_9 bias1 VCC VCC dummy_9
+ bias1 dummy_9 bias1 dummy_9 bias1 VCC dummy_9 bias1 VCC dummy_9 dummy_9 bias1 dummy_9
+ bias1 dummy_9 dummy_9 VCC VCC VCC dummy_9 bias1 VCC VCC VCC dummy_9 dummy_9 dummy_9
+ bias1 bias1 dummy_9 dummy_9 VCC VCC VCC bias1 bias1 dummy_9 dummy_9 VCC VCC dummy_9
+ dummy_9 dummy_9 VCC VCC VCC VCC bias1 VCC VCC dummy_9 bias1 dummy_9 dummy_9 dummy_9
+ bias1 bias1 dummy_9 dummy_9 dummy_9 dummy_9 bias1 dummy_9 VCC VCC dummy_9 bias1
+ dummy_9 dummy_9 bias1 dummy_9 dummy_9 VCC VCC dummy_9 dummy_9 VCC dummy_9 dummy_9
+ bias1 dummy_9 dummy_9 bias1 dummy_9 dummy_9 bias1 dummy_9 VCC bias1 dummy_9 bias1
+ VCC dummy_9 bias1 VCC dummy_9 dummy_9 dummy_9 VCC VCC dummy_9 bias1 VCC dummy_9
+ dummy_9 bias1 dummy_9 VCC dummy_9 dummy_9 dummy_9 VCC bias1 dummy_9 dummy_9 VCC
+ VCC dummy_9 bias1 dummy_9 bias1 dummy_9 dummy_9 dummy_9 dummy_9 dummy_9 VCC VCC
+ dummy_9 bias1 dummy_9 bias1 bias1 dummy_9 bias1 dummy_9 dummy_9 VCC VCC VCC dummy_9
+ dummy_9 dummy_9 bias1 dummy_9 dummy_9 dummy_9 bias1 VCC VCC bias1 dummy_9 dummy_9
+ dummy_9 VCC dummy_9 VCC VCC VSS dummy_9 dummy_9 sky130_fd_pr__pfet_01v8_E769TZ
XXM6_2 bias3 bias3 VSS VSS sky130_fd_pr__nfet_01v8_VT3ZQW
XXM8 VSS bias21 bias21 VSS sky130_fd_pr__nfet_01v8_VT3ZQW
XXM2_dummy_2 dummy_2 dummy_2 VB_A VB_A dummy_2 dummy_2 VB_A dummy_2 VCC VCC dummy_2
+ dummy_2 dummy_2 VB_A VCC dummy_2 dummy_2 VCC dummy_2 VCC VCC VB_A dummy_2 VCC VB_A
+ dummy_2 VCC dummy_2 VB_A VB_A dummy_2 VB_A dummy_2 dummy_2 dummy_2 dummy_2 dummy_2
+ VCC dummy_2 VCC VCC dummy_2 dummy_2 VCC dummy_2 dummy_2 dummy_2 VB_A VB_A VB_A VCC
+ dummy_2 VB_A VB_A VCC VB_A dummy_2 VCC VB_A dummy_2 VCC dummy_2 VB_A dummy_2 dummy_2
+ VCC dummy_2 dummy_2 VSS sky130_fd_pr__pfet_01v8_UDMRD5
Xsky130_fd_pr__pfet_01v8_RRU5GE_0 IB VCC m1_44990_37960# VCC VCC IB VCC IB VCC VCC
+ m1_44990_37960# m1_44990_37960# VSS sky130_fd_pr__pfet_01v8_RRU5GE
XXM6_3 bias3 bias3 VSS VSS sky130_fd_pr__nfet_01v8_VT3ZQW
XXM9 VCC VCC bias1 VCC bias1 VCC m9m10 bias1 VCC VCC m9m10 bias1 VCC VCC m9m10 VCC
+ m9m10 bias1 bias1 VCC VCC m9m10 bias1 VCC VCC VCC VCC bias1 VCC VCC m9m10 bias1
+ VCC m9m10 m9m10 VCC VCC VCC bias1 VCC bias1 VCC bias1 m9m10 VCC m9m10 bias1 VCC
+ m9m10 bias1 VCC VCC VCC m9m10 VCC VCC bias1 m9m10 m9m10 bias1 VCC VCC bias1 bias1
+ VCC VCC m9m10 VCC bias1 m9m10 bias1 m9m10 VCC m9m10 bias1 VCC VCC VCC m9m10 VCC
+ VCC VCC VCC VCC bias1 VCC bias1 m9m10 bias1 bias1 bias1 VCC m9m10 VCC bias1 VCC
+ m9m10 VCC m9m10 bias1 VCC VCC VCC VCC bias1 VCC VCC VCC m9m10 bias1 m9m10 VCC VCC
+ bias1 VCC bias1 m9m10 VCC VCC VCC VCC bias1 VCC m9m10 VCC m9m10 bias1 bias1 m9m10
+ m9m10 VCC VCC bias1 VCC VCC VCC bias1 VCC m9m10 m9m10 VCC VCC VCC VCC m9m10 VCC
+ VCC bias1 bias1 VCC VCC m9m10 VCC m9m10 m9m10 VCC VCC VCC m9m10 bias1 m9m10 VCC
+ bias1 VCC m9m10 VCC VCC VCC VCC m9m10 VCC m9m10 VCC VCC VCC bias1 VCC bias1 bias1
+ m9m10 bias1 VCC m9m10 bias1 VCC bias1 VCC VCC VCC VCC VCC bias1 bias1 m9m10 bias1
+ bias1 VCC bias1 m9m10 VCC VCC VCC bias1 bias1 VCC VCC VCC VCC bias1 m9m10 bias1
+ m9m10 m9m10 VCC m9m10 bias1 VCC VCC bias1 VCC bias1 VCC m9m10 m9m10 m9m10 bias1
+ VCC VCC m9m10 bias1 bias1 m9m10 m9m10 bias1 VCC m9m10 VCC bias1 VCC VCC m9m10 bias1
+ VCC bias1 m9m10 bias1 VCC m9m10 bias1 VCC m9m10 m9m10 bias1 m9m10 bias1 VCC VCC
+ VCC VCC VCC m9m10 bias1 VCC VCC VCC m9m10 m9m10 VCC bias1 bias1 m9m10 VCC VCC VCC
+ VCC bias1 bias1 m9m10 m9m10 VCC VCC VCC VCC VCC VCC VCC VCC VCC bias1 VCC VCC VCC
+ bias1 m9m10 m9m10 m9m10 bias1 bias1 m9m10 m9m10 VCC VCC bias1 VCC VCC VCC bias1
+ VCC m9m10 bias1 VCC VCC VCC VCC VCC m9m10 VCC VCC m9m10 bias1 VCC VCC bias1 VCC
+ m9m10 bias1 m9m10 VCC bias1 m9m10 bias1 VCC m9m10 bias1 VCC m9m10 m9m10 VCC VCC
+ VCC m9m10 bias1 VCC VCC m9m10 bias1 VCC VCC VCC VCC VCC VCC bias1 VCC m9m10 VCC
+ VCC m9m10 bias1 m9m10 bias1 VCC m9m10 VCC m9m10 VCC VCC VCC m9m10 bias1 m9m10 bias1
+ bias1 VCC bias1 m9m10 m9m10 VCC VCC VCC m9m10 m9m10 m9m10 bias1 m9m10 m9m10 VCC
+ bias1 VCC VCC bias1 m9m10 VCC VCC VCC VCC VCC VCC VSS m9m10 VCC sky130_fd_pr__pfet_01v8_F76D73
XXM2_dummy_3 VB_A dummy_2 VCC dummy_2 VSS sky130_fd_pr__pfet_01v8_SKU9VM
Xsky130_fd_pr__pfet_01v8_C2U9V5_0 IB dummy_100 VCC dummy_100 VSS sky130_fd_pr__pfet_01v8_C2U9V5
XXM2_dummy_4 VB_A dummy_2 VCC dummy_2 VSS sky130_fd_pr__pfet_01v8_SKU9VM
XXM2_dummy_5 VB_A dummy_2 VCC dummy_2 VSS sky130_fd_pr__pfet_01v8_SKU9VM
Xsky130_fd_pr__nfet_01v8_AH5E2K_0 dummy_3 dummy_3 VB_B VSS sky130_fd_pr__nfet_01v8_AH5E2K
XXM2_1 m1m2 VB_A bias1 m1m2 VB_A bias1 VCC VCC bias1 bias1 bias1 VB_A VCC bias1 VCC
+ m1m2 VCC VCC VB_A m1m2 VCC VB_A m1m2 m1m2 VB_A VB_A bias1 VB_A bias1 bias1 m1m2
+ bias1 VCC bias1 VCC VCC m1m2 m1m2 VCC m1m2 m1m2 m1m2 VB_A VB_A VB_A VCC bias1 VB_A
+ VCC VB_A bias1 VCC VB_A bias1 VCC VB_A bias1 m1m2 m1m2 m1m2 VSS sky130_fd_pr__pfet_01v8_UDM5A5
XXM2_dummy_6 VB_A dummy_2 VCC dummy_2 VSS sky130_fd_pr__pfet_01v8_SKU9VM
Xsky130_fd_pr__nfet_01v8_3ZAA45_0 m11m12 VSS bias21 VSS sky130_fd_pr__nfet_01v8_3ZAA45
XXM3_dummy_10 dummy_3 dummy_3 VB_B VSS sky130_fd_pr__nfet_01v8_AH5E2K
Xsky130_fd_pr__nfet_01v8_MHE452_0 dummy_4 bias3 dummy_4 dummy_4 bias3 dummy_4 bias3
+ dummy_4 bias3 dummy_4 dummy_4 dummy_4 dummy_4 dummy_4 bias3 dummy_4 dummy_4 bias3
+ VSS sky130_fd_pr__nfet_01v8_MHE452
XXM2_dummy_7 VB_A dummy_2 VCC dummy_2 VSS sky130_fd_pr__pfet_01v8_SKU9VM
Xsky130_fd_pr__pfet_01v8_F76D73_0 m1m2 m1m2 bias1 VCC bias1 m1m2 VCC bias1 VCC VCC
+ VCC bias1 m1m2 VCC VCC m1m2 VCC bias1 bias1 VCC VCC VCC bias1 m1m2 m1m2 m1m2 m1m2
+ bias1 VCC m1m2 VCC bias1 VCC VCC VCC m1m2 m1m2 VCC bias1 VCC bias1 m1m2 bias1 VCC
+ m1m2 VCC bias1 m1m2 VCC bias1 m1m2 VCC VCC VCC VCC VCC bias1 VCC VCC bias1 m1m2
+ m1m2 bias1 bias1 VCC VCC VCC m1m2 bias1 VCC bias1 VCC m1m2 VCC bias1 m1m2 VCC VCC
+ VCC VCC VCC m1m2 VCC m1m2 bias1 m1m2 bias1 VCC bias1 bias1 bias1 VCC VCC VCC bias1
+ m1m2 VCC m1m2 VCC bias1 m1m2 m1m2 VCC VCC bias1 VCC m1m2 m1m2 VCC bias1 VCC m1m2
+ m1m2 bias1 VCC bias1 VCC VCC m1m2 m1m2 VCC bias1 VCC VCC m1m2 VCC bias1 bias1 VCC
+ VCC m1m2 VCC bias1 m1m2 VCC m1m2 bias1 VCC VCC VCC m1m2 m1m2 VCC VCC VCC VCC VCC
+ bias1 bias1 m1m2 m1m2 VCC m1m2 VCC VCC m1m2 VCC VCC VCC bias1 VCC m1m2 bias1 VCC
+ VCC m1m2 m1m2 m1m2 VCC VCC m1m2 VCC VCC VCC m1m2 bias1 m1m2 bias1 bias1 VCC bias1
+ VCC VCC bias1 VCC bias1 VCC m1m2 VCC m1m2 m1m2 bias1 bias1 VCC bias1 bias1 VCC bias1
+ VCC m1m2 m1m2 VCC bias1 bias1 VCC VCC m1m2 m1m2 bias1 VCC bias1 VCC VCC VCC VCC
+ bias1 m1m2 m1m2 bias1 m1m2 bias1 VCC VCC VCC VCC bias1 m1m2 m1m2 VCC bias1 bias1
+ VCC VCC bias1 VCC VCC m1m2 bias1 VCC VCC VCC bias1 m1m2 bias1 VCC bias1 VCC VCC
+ bias1 VCC VCC VCC bias1 VCC bias1 m1m2 m1m2 VCC VCC VCC VCC bias1 VCC VCC VCC VCC
+ VCC m1m2 bias1 bias1 VCC m1m2 VCC VCC VCC bias1 bias1 VCC VCC VCC VCC m1m2 m1m2
+ m1m2 VCC VCC VCC VCC bias1 VCC VCC m1m2 bias1 VCC VCC VCC bias1 bias1 VCC VCC m1m2
+ m1m2 bias1 m1m2 VCC VCC bias1 m1m2 VCC bias1 m1m2 m1m2 VCC VCC m1m2 VCC VCC m1m2
+ VCC bias1 m1m2 m1m2 bias1 m1m2 VCC bias1 VCC VCC bias1 VCC bias1 VCC VCC bias1 VCC
+ VCC VCC m1m2 VCC VCC VCC bias1 VCC m1m2 VCC bias1 m1m2 VCC m1m2 m1m2 m1m2 VCC bias1
+ m1m2 VCC VCC VCC VCC bias1 VCC bias1 m1m2 VCC m1m2 VCC m1m2 VCC VCC VCC bias1 VCC
+ bias1 bias1 m1m2 bias1 VCC VCC VCC VCC VCC VCC VCC VCC bias1 VCC VCC m1m2 bias1
+ VCC VCC bias1 VCC m1m2 m1m2 VCC m1m2 VCC VCC VSS VCC m1m2 sky130_fd_pr__pfet_01v8_F76D73
Xsky130_fd_pr__pfet_01v8_UDM5A5_0 m9m10 VB_A OUT m9m10 VB_A OUT VCC VCC OUT OUT OUT
+ VB_A VCC OUT VCC m9m10 VCC VCC VB_A m9m10 VCC VB_A m9m10 m9m10 VB_A VB_A OUT VB_A
+ OUT OUT m9m10 OUT VCC OUT VCC VCC m9m10 m9m10 VCC m9m10 m9m10 m9m10 VB_A VB_A VB_A
+ VCC OUT VB_A VCC VB_A OUT VCC VB_A OUT VCC VB_A OUT m9m10 m9m10 m9m10 VSS sky130_fd_pr__pfet_01v8_UDM5A5
XXM9_dummy_1 dummy_9 dummy_9 bias1 VCC bias1 dummy_9 dummy_9 bias1 VCC VCC dummy_9
+ bias1 dummy_9 VCC VCC dummy_9 dummy_9 dummy_9 bias1 bias1 VCC VCC dummy_9 bias1
+ dummy_9 dummy_9 dummy_9 dummy_9 bias1 VCC dummy_9 dummy_9 bias1 VCC dummy_9 dummy_9
+ dummy_9 dummy_9 VCC bias1 VCC bias1 dummy_9 bias1 dummy_9 dummy_9 dummy_9 bias1
+ dummy_9 dummy_9 bias1 dummy_9 bias1 VCC VCC dummy_9 VCC VCC bias1 dummy_9 dummy_9
+ bias1 dummy_9 dummy_9 bias1 bias1 VCC VCC dummy_9 dummy_9 bias1 dummy_9 bias1 dummy_9
+ dummy_9 dummy_9 bias1 dummy_9 VCC VCC dummy_9 VCC VCC dummy_9 VCC dummy_9 bias1
+ dummy_9 bias1 dummy_9 bias1 bias1 bias1 VCC dummy_9 VCC bias1 dummy_9 dummy_9 dummy_9
+ dummy_9 bias1 dummy_9 dummy_9 VCC bias1 VCC VCC dummy_9 dummy_9 dummy_9 bias1 dummy_9
+ dummy_9 dummy_9 bias1 VCC bias1 dummy_9 VCC dummy_9 dummy_9 dummy_9 VCC bias1 VCC
+ dummy_9 dummy_9 dummy_9 bias1 bias1 dummy_9 dummy_9 dummy_9 dummy_9 VCC bias1 dummy_9
+ VCC dummy_9 bias1 VCC dummy_9 VCC dummy_9 dummy_9 dummy_9 VCC VCC dummy_9 VCC VCC
+ bias1 bias1 dummy_9 dummy_9 dummy_9 dummy_9 dummy_9 dummy_9 dummy_9 VCC VCC dummy_9
+ dummy_9 bias1 dummy_9 dummy_9 bias1 VCC dummy_9 dummy_9 dummy_9 dummy_9 VCC dummy_9
+ dummy_9 dummy_9 VCC VCC dummy_9 bias1 dummy_9 bias1 bias1 dummy_9 bias1 VCC dummy_9
+ bias1 VCC bias1 VCC dummy_9 VCC dummy_9 dummy_9 bias1 bias1 dummy_9 bias1 bias1
+ VCC bias1 dummy_9 dummy_9 dummy_9 VCC bias1 bias1 VCC VCC dummy_9 dummy_9 bias1
+ dummy_9 bias1 dummy_9 dummy_9 VCC bias1 dummy_9 bias1 dummy_9 dummy_9 bias1 dummy_9
+ bias1 VCC dummy_9 dummy_9 dummy_9 bias1 dummy_9 dummy_9 dummy_9 bias1 bias1 dummy_9
+ dummy_9 bias1 VCC dummy_9 dummy_9 bias1 VCC VCC dummy_9 bias1 dummy_9 bias1 dummy_9
+ bias1 VCC dummy_9 bias1 VCC dummy_9 dummy_9 bias1 dummy_9 bias1 dummy_9 dummy_9
+ VCC VCC VCC dummy_9 bias1 VCC VCC VCC dummy_9 dummy_9 dummy_9 bias1 bias1 dummy_9
+ dummy_9 VCC VCC VCC bias1 bias1 dummy_9 dummy_9 VCC VCC dummy_9 dummy_9 dummy_9
+ VCC VCC VCC VCC bias1 VCC VCC dummy_9 bias1 dummy_9 dummy_9 dummy_9 bias1 bias1
+ dummy_9 dummy_9 dummy_9 dummy_9 bias1 dummy_9 VCC VCC dummy_9 bias1 dummy_9 dummy_9
+ bias1 dummy_9 dummy_9 VCC VCC dummy_9 dummy_9 VCC dummy_9 dummy_9 bias1 dummy_9
+ dummy_9 bias1 dummy_9 dummy_9 bias1 dummy_9 VCC bias1 dummy_9 bias1 VCC dummy_9
+ bias1 VCC dummy_9 dummy_9 dummy_9 VCC VCC dummy_9 bias1 VCC dummy_9 dummy_9 bias1
+ dummy_9 VCC dummy_9 dummy_9 dummy_9 VCC bias1 dummy_9 dummy_9 VCC VCC dummy_9 bias1
+ dummy_9 bias1 dummy_9 dummy_9 dummy_9 dummy_9 dummy_9 VCC VCC dummy_9 bias1 dummy_9
+ bias1 bias1 dummy_9 bias1 dummy_9 dummy_9 VCC VCC VCC dummy_9 dummy_9 dummy_9 bias1
+ dummy_9 dummy_9 dummy_9 bias1 VCC VCC bias1 dummy_9 dummy_9 dummy_9 VCC dummy_9
+ VCC VCC VSS dummy_9 dummy_9 sky130_fd_pr__pfet_01v8_E769TZ
XXM2_dummy_9 VB_A dummy_2 VCC dummy_2 VSS sky130_fd_pr__pfet_01v8_SKU9VM
XXM5_dummy_1 VCC IN_P IN_P dummy_5 IN_P VCC dummy_5 VCC dummy_5 dummy_5 dummy_5 dummy_5
+ IN_P dummy_5 dummy_5 VCC dummy_5 IN_P dummy_5 dummy_5 VCC dummy_5 IN_P IN_P dummy_5
+ VCC IN_P IN_P IN_P VCC VCC dummy_5 VCC IN_P IN_P VCC IN_P dummy_5 dummy_5 dummy_5
+ dummy_5 IN_P VCC dummy_5 dummy_5 dummy_5 dummy_5 IN_P VCC dummy_5 dummy_5 VCC dummy_5
+ dummy_5 VCC VCC dummy_5 dummy_5 dummy_5 dummy_5 dummy_5 dummy_5 dummy_5 VCC IN_P
+ dummy_5 IN_P VCC VSS sky130_fd_pr__pfet_01v8_8DHNHY
XXM9_dummy_3 VCC bias1 dummy_9 dummy_9 VSS sky130_fd_pr__pfet_01v8_SLZ774
XXM5_dummy_3 dummy_5 IN_P VCC dummy_5 VSS sky130_fd_pr__pfet_01v8_MGA63L
XXM9_dummy_4 VCC bias1 dummy_9 dummy_9 VSS sky130_fd_pr__pfet_01v8_ZLZ7XS
XXM5_dummy_4 dummy_5 IN_P VCC dummy_5 VSS sky130_fd_pr__pfet_01v8_MGA63L
Xsky130_fd_pr__pfet_01v8_UDMRD5_0 dummy_2 dummy_2 VB_A VB_A dummy_2 dummy_2 VB_A dummy_2
+ VCC VCC dummy_2 dummy_2 dummy_2 VB_A VCC dummy_2 dummy_2 VCC dummy_2 VCC VCC VB_A
+ dummy_2 VCC VB_A dummy_2 VCC dummy_2 VB_A VB_A dummy_2 VB_A dummy_2 dummy_2 dummy_2
+ dummy_2 dummy_2 VCC dummy_2 VCC VCC dummy_2 dummy_2 VCC dummy_2 dummy_2 dummy_2
+ VB_A VB_A VB_A VCC dummy_2 VB_A VB_A VCC VB_A dummy_2 VCC VB_A dummy_2 VCC dummy_2
+ VB_A dummy_2 dummy_2 VCC dummy_2 dummy_2 VSS sky130_fd_pr__pfet_01v8_UDMRD5
XXM9_dummy_5 VCC bias1 dummy_9 dummy_9 VSS sky130_fd_pr__pfet_01v8_ZLZ7XS
XXM9_1 VCC VCC bias1 VCC bias1 VCC m9m10 bias1 VCC VCC m9m10 bias1 VCC VCC m9m10 VCC
+ m9m10 bias1 bias1 VCC VCC m9m10 bias1 VCC VCC VCC VCC bias1 VCC VCC m9m10 bias1
+ VCC m9m10 m9m10 VCC VCC VCC bias1 VCC bias1 VCC bias1 m9m10 VCC m9m10 bias1 VCC
+ m9m10 bias1 VCC VCC VCC m9m10 VCC VCC bias1 m9m10 m9m10 bias1 VCC VCC bias1 bias1
+ VCC VCC m9m10 VCC bias1 m9m10 bias1 m9m10 VCC m9m10 bias1 VCC VCC VCC m9m10 VCC
+ VCC VCC VCC VCC bias1 VCC bias1 m9m10 bias1 bias1 bias1 VCC m9m10 VCC bias1 VCC
+ m9m10 VCC m9m10 bias1 VCC VCC VCC VCC bias1 VCC VCC VCC m9m10 bias1 m9m10 VCC VCC
+ bias1 VCC bias1 m9m10 VCC VCC VCC VCC bias1 VCC m9m10 VCC m9m10 bias1 bias1 m9m10
+ m9m10 VCC VCC bias1 VCC VCC VCC bias1 VCC m9m10 m9m10 VCC VCC VCC VCC m9m10 VCC
+ VCC bias1 bias1 VCC VCC m9m10 VCC m9m10 m9m10 VCC VCC VCC m9m10 bias1 m9m10 VCC
+ bias1 VCC m9m10 VCC VCC VCC VCC m9m10 VCC m9m10 VCC VCC VCC bias1 VCC bias1 bias1
+ m9m10 bias1 VCC m9m10 bias1 VCC bias1 VCC VCC VCC VCC VCC bias1 bias1 m9m10 bias1
+ bias1 VCC bias1 m9m10 VCC VCC VCC bias1 bias1 VCC VCC VCC VCC bias1 m9m10 bias1
+ m9m10 m9m10 VCC m9m10 bias1 VCC VCC bias1 VCC bias1 VCC m9m10 m9m10 m9m10 bias1
+ VCC VCC m9m10 bias1 bias1 m9m10 m9m10 bias1 VCC m9m10 VCC bias1 VCC VCC m9m10 bias1
+ VCC bias1 m9m10 bias1 VCC m9m10 bias1 VCC m9m10 m9m10 bias1 m9m10 bias1 VCC VCC
+ VCC VCC VCC m9m10 bias1 VCC VCC VCC m9m10 m9m10 VCC bias1 bias1 m9m10 VCC VCC VCC
+ VCC bias1 bias1 m9m10 m9m10 VCC VCC VCC VCC VCC VCC VCC VCC VCC bias1 VCC VCC VCC
+ bias1 m9m10 m9m10 m9m10 bias1 bias1 m9m10 m9m10 VCC VCC bias1 VCC VCC VCC bias1
+ VCC m9m10 bias1 VCC VCC VCC VCC VCC m9m10 VCC VCC m9m10 bias1 VCC VCC bias1 VCC
+ m9m10 bias1 m9m10 VCC bias1 m9m10 bias1 VCC m9m10 bias1 VCC m9m10 m9m10 VCC VCC
+ VCC m9m10 bias1 VCC VCC m9m10 bias1 VCC VCC VCC VCC VCC VCC bias1 VCC m9m10 VCC
+ VCC m9m10 bias1 m9m10 bias1 VCC m9m10 VCC m9m10 VCC VCC VCC m9m10 bias1 m9m10 bias1
+ bias1 VCC bias1 m9m10 m9m10 VCC VCC VCC m9m10 m9m10 m9m10 bias1 m9m10 m9m10 VCC
+ bias1 VCC VCC bias1 m9m10 VCC VCC VCC VCC VCC VCC VSS m9m10 VCC sky130_fd_pr__pfet_01v8_F76D73
XXM9_dummy_20 VCC bias1 dummy_9 dummy_9 VSS sky130_fd_pr__pfet_01v8_ZLZ7XS
XXM5_dummy_5 dummy_5 IN_P VCC dummy_5 VSS sky130_fd_pr__pfet_01v8_MGA63L
XXM9_dummy_6 VCC bias1 dummy_9 dummy_9 VSS sky130_fd_pr__pfet_01v8_ZLZ7XS
XXM9_dummy_10 VCC bias1 dummy_9 dummy_9 VSS sky130_fd_pr__pfet_01v8_ZLZ7XS
XXM9_2 VCC VCC bias1 VCC bias1 VCC m9m10 bias1 VCC VCC m9m10 bias1 VCC VCC m9m10 VCC
+ m9m10 bias1 bias1 VCC VCC m9m10 bias1 VCC VCC VCC VCC bias1 VCC VCC m9m10 bias1
+ VCC m9m10 m9m10 VCC VCC VCC bias1 VCC bias1 VCC bias1 m9m10 VCC m9m10 bias1 VCC
+ m9m10 bias1 VCC VCC VCC m9m10 VCC VCC bias1 m9m10 m9m10 bias1 VCC VCC bias1 bias1
+ VCC VCC m9m10 VCC bias1 m9m10 bias1 m9m10 VCC m9m10 bias1 VCC VCC VCC m9m10 VCC
+ VCC VCC VCC VCC bias1 VCC bias1 m9m10 bias1 bias1 bias1 VCC m9m10 VCC bias1 VCC
+ m9m10 VCC m9m10 bias1 VCC VCC VCC VCC bias1 VCC VCC VCC m9m10 bias1 m9m10 VCC VCC
+ bias1 VCC bias1 m9m10 VCC VCC VCC VCC bias1 VCC m9m10 VCC m9m10 bias1 bias1 m9m10
+ m9m10 VCC VCC bias1 VCC VCC VCC bias1 VCC m9m10 m9m10 VCC VCC VCC VCC m9m10 VCC
+ VCC bias1 bias1 VCC VCC m9m10 VCC m9m10 m9m10 VCC VCC VCC m9m10 bias1 m9m10 VCC
+ bias1 VCC m9m10 VCC VCC VCC VCC m9m10 VCC m9m10 VCC VCC VCC bias1 VCC bias1 bias1
+ m9m10 bias1 VCC m9m10 bias1 VCC bias1 VCC VCC VCC VCC VCC bias1 bias1 m9m10 bias1
+ bias1 VCC bias1 m9m10 VCC VCC VCC bias1 bias1 VCC VCC VCC VCC bias1 m9m10 bias1
+ m9m10 m9m10 VCC m9m10 bias1 VCC VCC bias1 VCC bias1 VCC m9m10 m9m10 m9m10 bias1
+ VCC VCC m9m10 bias1 bias1 m9m10 m9m10 bias1 VCC m9m10 VCC bias1 VCC VCC m9m10 bias1
+ VCC bias1 m9m10 bias1 VCC m9m10 bias1 VCC m9m10 m9m10 bias1 m9m10 bias1 VCC VCC
+ VCC VCC VCC m9m10 bias1 VCC VCC VCC m9m10 m9m10 VCC bias1 bias1 m9m10 VCC VCC VCC
+ VCC bias1 bias1 m9m10 m9m10 VCC VCC VCC VCC VCC VCC VCC VCC VCC bias1 VCC VCC VCC
+ bias1 m9m10 m9m10 m9m10 bias1 bias1 m9m10 m9m10 VCC VCC bias1 VCC VCC VCC bias1
+ VCC m9m10 bias1 VCC VCC VCC VCC VCC m9m10 VCC VCC m9m10 bias1 VCC VCC bias1 VCC
+ m9m10 bias1 m9m10 VCC bias1 m9m10 bias1 VCC m9m10 bias1 VCC m9m10 m9m10 VCC VCC
+ VCC m9m10 bias1 VCC VCC m9m10 bias1 VCC VCC VCC VCC VCC VCC bias1 VCC m9m10 VCC
+ VCC m9m10 bias1 m9m10 bias1 VCC m9m10 VCC m9m10 VCC VCC VCC m9m10 bias1 m9m10 bias1
+ bias1 VCC bias1 m9m10 m9m10 VCC VCC VCC m9m10 m9m10 m9m10 bias1 m9m10 m9m10 VCC
+ bias1 VCC VCC bias1 m9m10 VCC VCC VCC VCC VCC VCC VSS m9m10 VCC sky130_fd_pr__pfet_01v8_F76D73
XXM5_dummy_6 dummy_5 IN_P VCC dummy_5 VSS sky130_fd_pr__pfet_01v8_MGA63L
XXM9_dummy_7 VCC bias1 dummy_9 dummy_9 VSS sky130_fd_pr__pfet_01v8_ZLZ7XS
XXM9_dummy_22 VCC bias1 dummy_9 dummy_9 VSS sky130_fd_pr__pfet_01v8_ZLZ7XS
XXM9_dummy_11 VCC bias1 dummy_9 dummy_9 VSS sky130_fd_pr__pfet_01v8_ZLZ7XS
XXM9_3 VCC VCC bias1 VCC bias1 VCC m9m10 bias1 VCC VCC m9m10 bias1 VCC VCC m9m10 VCC
+ m9m10 bias1 bias1 VCC VCC m9m10 bias1 VCC VCC VCC VCC bias1 VCC VCC m9m10 bias1
+ VCC m9m10 m9m10 VCC VCC VCC bias1 VCC bias1 VCC bias1 m9m10 VCC m9m10 bias1 VCC
+ m9m10 bias1 VCC VCC VCC m9m10 VCC VCC bias1 m9m10 m9m10 bias1 VCC VCC bias1 bias1
+ VCC VCC m9m10 VCC bias1 m9m10 bias1 m9m10 VCC m9m10 bias1 VCC VCC VCC m9m10 VCC
+ VCC VCC VCC VCC bias1 VCC bias1 m9m10 bias1 bias1 bias1 VCC m9m10 VCC bias1 VCC
+ m9m10 VCC m9m10 bias1 VCC VCC VCC VCC bias1 VCC VCC VCC m9m10 bias1 m9m10 VCC VCC
+ bias1 VCC bias1 m9m10 VCC VCC VCC VCC bias1 VCC m9m10 VCC m9m10 bias1 bias1 m9m10
+ m9m10 VCC VCC bias1 VCC VCC VCC bias1 VCC m9m10 m9m10 VCC VCC VCC VCC m9m10 VCC
+ VCC bias1 bias1 VCC VCC m9m10 VCC m9m10 m9m10 VCC VCC VCC m9m10 bias1 m9m10 VCC
+ bias1 VCC m9m10 VCC VCC VCC VCC m9m10 VCC m9m10 VCC VCC VCC bias1 VCC bias1 bias1
+ m9m10 bias1 VCC m9m10 bias1 VCC bias1 VCC VCC VCC VCC VCC bias1 bias1 m9m10 bias1
+ bias1 VCC bias1 m9m10 VCC VCC VCC bias1 bias1 VCC VCC VCC VCC bias1 m9m10 bias1
+ m9m10 m9m10 VCC m9m10 bias1 VCC VCC bias1 VCC bias1 VCC m9m10 m9m10 m9m10 bias1
+ VCC VCC m9m10 bias1 bias1 m9m10 m9m10 bias1 VCC m9m10 VCC bias1 VCC VCC m9m10 bias1
+ VCC bias1 m9m10 bias1 VCC m9m10 bias1 VCC m9m10 m9m10 bias1 m9m10 bias1 VCC VCC
+ VCC VCC VCC m9m10 bias1 VCC VCC VCC m9m10 m9m10 VCC bias1 bias1 m9m10 VCC VCC VCC
+ VCC bias1 bias1 m9m10 m9m10 VCC VCC VCC VCC VCC VCC VCC VCC VCC bias1 VCC VCC VCC
+ bias1 m9m10 m9m10 m9m10 bias1 bias1 m9m10 m9m10 VCC VCC bias1 VCC VCC VCC bias1
+ VCC m9m10 bias1 VCC VCC VCC VCC VCC m9m10 VCC VCC m9m10 bias1 VCC VCC bias1 VCC
+ m9m10 bias1 m9m10 VCC bias1 m9m10 bias1 VCC m9m10 bias1 VCC m9m10 m9m10 VCC VCC
+ VCC m9m10 bias1 VCC VCC m9m10 bias1 VCC VCC VCC VCC VCC VCC bias1 VCC m9m10 VCC
+ VCC m9m10 bias1 m9m10 bias1 VCC m9m10 VCC m9m10 VCC VCC VCC m9m10 bias1 m9m10 bias1
+ bias1 VCC bias1 m9m10 m9m10 VCC VCC VCC m9m10 m9m10 m9m10 bias1 m9m10 m9m10 VCC
+ bias1 VCC VCC bias1 m9m10 VCC VCC VCC VCC VCC VCC VSS m9m10 VCC sky130_fd_pr__pfet_01v8_F76D73
XXM11_1 OUT OUT VB_B OUT VB_B VB_B VB_B VB_B m11m12 m11m12 m11m12 m11m12 OUT OUT VB_B
+ OUT OUT VB_B OUT OUT m11m12 VB_B m11m12 m11m12 m11m12 m11m12 m11m12 VB_B VB_B OUT
+ OUT VB_B OUT VB_B OUT VB_B VB_B m11m12 VB_B m11m12 m11m12 m11m12 m11m12 OUT OUT
+ VSS sky130_fd_pr__nfet_01v8_QP5WRD
XXM5_dummy_7 dummy_5 IN_P VCC dummy_5 VSS sky130_fd_pr__pfet_01v8_MGA63L
XXM9_dummy_8 VCC bias1 dummy_9 dummy_9 VSS sky130_fd_pr__pfet_01v8_ZLZ7XS
Xsky130_fd_pr__nfet_01v8_SCE452_0 dummy_4 bias3 dummy_4 VSS sky130_fd_pr__nfet_01v8_SCE452
XXM9_4 VCC VCC bias1 VCC bias1 VCC m9m10 bias1 VCC VCC m9m10 bias1 VCC VCC m9m10 VCC
+ m9m10 bias1 bias1 VCC VCC m9m10 bias1 VCC VCC VCC VCC bias1 VCC VCC m9m10 bias1
+ VCC m9m10 m9m10 VCC VCC VCC bias1 VCC bias1 VCC bias1 m9m10 VCC m9m10 bias1 VCC
+ m9m10 bias1 VCC VCC VCC m9m10 VCC VCC bias1 m9m10 m9m10 bias1 VCC VCC bias1 bias1
+ VCC VCC m9m10 VCC bias1 m9m10 bias1 m9m10 VCC m9m10 bias1 VCC VCC VCC m9m10 VCC
+ VCC VCC VCC VCC bias1 VCC bias1 m9m10 bias1 bias1 bias1 VCC m9m10 VCC bias1 VCC
+ m9m10 VCC m9m10 bias1 VCC VCC VCC VCC bias1 VCC VCC VCC m9m10 bias1 m9m10 VCC VCC
+ bias1 VCC bias1 m9m10 VCC VCC VCC VCC bias1 VCC m9m10 VCC m9m10 bias1 bias1 m9m10
+ m9m10 VCC VCC bias1 VCC VCC VCC bias1 VCC m9m10 m9m10 VCC VCC VCC VCC m9m10 VCC
+ VCC bias1 bias1 VCC VCC m9m10 VCC m9m10 m9m10 VCC VCC VCC m9m10 bias1 m9m10 VCC
+ bias1 VCC m9m10 VCC VCC VCC VCC m9m10 VCC m9m10 VCC VCC VCC bias1 VCC bias1 bias1
+ m9m10 bias1 VCC m9m10 bias1 VCC bias1 VCC VCC VCC VCC VCC bias1 bias1 m9m10 bias1
+ bias1 VCC bias1 m9m10 VCC VCC VCC bias1 bias1 VCC VCC VCC VCC bias1 m9m10 bias1
+ m9m10 m9m10 VCC m9m10 bias1 VCC VCC bias1 VCC bias1 VCC m9m10 m9m10 m9m10 bias1
+ VCC VCC m9m10 bias1 bias1 m9m10 m9m10 bias1 VCC m9m10 VCC bias1 VCC VCC m9m10 bias1
+ VCC bias1 m9m10 bias1 VCC m9m10 bias1 VCC m9m10 m9m10 bias1 m9m10 bias1 VCC VCC
+ VCC VCC VCC m9m10 bias1 VCC VCC VCC m9m10 m9m10 VCC bias1 bias1 m9m10 VCC VCC VCC
+ VCC bias1 bias1 m9m10 m9m10 VCC VCC VCC VCC VCC VCC VCC VCC VCC bias1 VCC VCC VCC
+ bias1 m9m10 m9m10 m9m10 bias1 bias1 m9m10 m9m10 VCC VCC bias1 VCC VCC VCC bias1
+ VCC m9m10 bias1 VCC VCC VCC VCC VCC m9m10 VCC VCC m9m10 bias1 VCC VCC bias1 VCC
+ m9m10 bias1 m9m10 VCC bias1 m9m10 bias1 VCC m9m10 bias1 VCC m9m10 m9m10 VCC VCC
+ VCC m9m10 bias1 VCC VCC m9m10 bias1 VCC VCC VCC VCC VCC VCC bias1 VCC m9m10 VCC
+ VCC m9m10 bias1 m9m10 bias1 VCC m9m10 VCC m9m10 VCC VCC VCC m9m10 bias1 m9m10 bias1
+ bias1 VCC bias1 m9m10 m9m10 VCC VCC VCC m9m10 m9m10 m9m10 bias1 m9m10 m9m10 VCC
+ bias1 VCC VCC bias1 m9m10 VCC VCC VCC VCC VCC VCC VSS m9m10 VCC sky130_fd_pr__pfet_01v8_F76D73
XXM9_dummy_12 VCC bias1 dummy_9 dummy_9 VSS sky130_fd_pr__pfet_01v8_ZLZ7XS
XXM5_dummy_8 dummy_5 IN_P VCC dummy_5 VSS sky130_fd_pr__pfet_01v8_MGA63L
XXM9_dummy_9 VCC bias1 dummy_9 dummy_9 VSS sky130_fd_pr__pfet_01v8_ZLZ7XS
XXM10 OUT VB_A m9m10 OUT VB_A m9m10 VCC VCC m9m10 m9m10 m9m10 VB_A VCC m9m10 VCC OUT
+ VCC VCC VB_A OUT VCC VB_A OUT OUT VB_A VB_A m9m10 VB_A m9m10 m9m10 OUT m9m10 VCC
+ m9m10 VCC VCC OUT OUT VCC OUT OUT OUT VB_A VB_A VB_A VCC m9m10 VB_A VCC VB_A m9m10
+ VCC VB_A m9m10 VCC VB_A m9m10 OUT OUT OUT VSS sky130_fd_pr__pfet_01v8_UDM5A5
Xsky130_fd_pr__nfet_01v8_SCE452_1 dummy_4 bias3 dummy_4 VSS sky130_fd_pr__nfet_01v8_SCE452
Xsky130_fd_pr__pfet_01v8_7DHACV_0 VCC IN_P IN_P m1_44990_37960# VCC VCC bias21 bias21
+ bias21 m1_44990_37960# IN_P m1_44990_37960# bias21 m1_44990_37960# IN_P bias21 m1_44990_37960#
+ VCC IN_P IN_P m1_44990_37960# VCC IN_P IN_P IN_P VCC VCC VCC IN_P IN_P IN_P bias21
+ bias21 bias21 m1_44990_37960# IN_P VCC m1_44990_37960# bias21 m1_44990_37960# bias21
+ IN_P VCC m1_44990_37960# bias21 VCC m1_44990_37960# VCC VCC bias21 m1_44990_37960#
+ bias21 m1_44990_37960# m1_44990_37960# bias21 m1_44990_37960# VCC bias21 IN_P VCC
+ VSS sky130_fd_pr__pfet_01v8_7DHACV
XXM9_dummy_13 VCC bias1 dummy_9 dummy_9 VSS sky130_fd_pr__pfet_01v8_ZLZ7XS
XXM100_1 IB VCC VCC m1_44990_37960# VCC IB m1_44990_37960# IB VCC m1_44990_37960#
+ VCC VCC VSS sky130_fd_pr__pfet_01v8_RRU5GE
XXM2_dummy_10 VB_A dummy_2 VCC dummy_2 VSS sky130_fd_pr__pfet_01v8_SKU9VM
XXM11 m11m12 m11m12 VB_B m11m12 VB_B VB_B VB_B VB_B OUT OUT OUT OUT m11m12 m11m12
+ VB_B m11m12 m11m12 VB_B m11m12 m11m12 OUT VB_B OUT OUT OUT OUT OUT VB_B VB_B m11m12
+ m11m12 VB_B m11m12 VB_B m11m12 VB_B VB_B OUT VB_B OUT OUT OUT OUT m11m12 m11m12
+ VSS sky130_fd_pr__nfet_01v8_QP5WRD
Xsky130_fd_pr__nfet_01v8_SCE452_2 dummy_4 bias3 dummy_4 VSS sky130_fd_pr__nfet_01v8_SCE452
Xsky130_fd_pr__nfet_01v8_WK8VRD_0 VB_B dummy_3 dummy_3 dummy_3 VB_B dummy_3 VB_B VB_B
+ VB_B VB_B dummy_3 dummy_3 dummy_3 dummy_3 dummy_3 dummy_3 VB_B dummy_3 dummy_3 dummy_3
+ VB_B dummy_3 dummy_3 dummy_3 VB_B dummy_3 dummy_3 dummy_3 dummy_3 VB_B dummy_3 dummy_3
+ VB_B VB_B dummy_3 dummy_3 VB_B dummy_3 VB_B dummy_3 VB_B VB_B dummy_3 VB_B dummy_3
+ dummy_3 dummy_3 dummy_3 dummy_3 dummy_3 dummy_3 VSS sky130_fd_pr__nfet_01v8_WK8VRD
XXM9_dummy_14 VCC bias1 dummy_9 dummy_9 VSS sky130_fd_pr__pfet_01v8_ZLZ7XS
C0 m9m10 OUT -1.25f
C1 bias21 VB_B 1.02f
C2 dummy_2 bias1 2.5f
C3 m1_44990_37960# IB 7.64f
C4 VCC OUT 13.6f
C5 dummy_2 bias21 0.891f
C6 dummy_5 bias21 0.398f
C7 VB_B dummy_3 33.2f
C8 VB_A dummy_2 33f
C9 IN_P dummy_5 31.3f
C10 IN_P IN_M 3.32f
C11 m3m4 VB_B 6.64f
C12 VCC dummy_100 8.42f
C13 bias1 OUT 1.55f
C14 OUT bias21 0.978f
C15 dummy_4 bias3 8.54f
C16 m11m12 VB_B 6.51f
C17 VB_A OUT 6.54f
C18 VCC bias3 42.5f
C19 OUT dummy_3 2.64f
C20 OUT m3m4 18.9f
C21 m9m10 VCC 0.147p
C22 bias21 bias3 10.1f
C23 m11m12 OUT -1.26f
C24 m9m10 bias1 80.7f
C25 VB_A bias3 0.977f
C26 bias21 dummy_4 0.403f
C27 IN_P bias3 0.727f
C28 dummy_5 m1_44990_37960# 15.5f
C29 IN_M m1_44990_37960# 10.4f
C30 bias1 VCC 0.849p
C31 VCC bias21 39.6f
C32 VB_A m9m10 5.59f
C33 dummy_9 m1m2 35f
C34 m3m4 bias3 1.29f
C35 VB_A VCC 37.3f
C36 VCC IN_P 29.6f
C37 dummy_4 m3m4 1.44f
C38 dummy_2 m1m2 2.66f
C39 m11m12 bias3 0.374f
C40 VB_A bias1 7.09f
C41 m11m12 dummy_4 1.08f
C42 m1_44990_37960# dummy_100 5.9f
C43 IB dummy_100 15.6f
C44 VB_A bias21 1.01f
C45 IN_P bias21 11.1f
C46 bias1 dummy_3 2.66f
C47 OUT m1m2 0.00992f
C48 bias21 dummy_3 0.965f
C49 bias1 m3m4 -1.25f
C50 bias21 m3m4 0.0154f
C51 m1_44990_37960# bias3 0.988f
C52 bias3 IB 0.619f
C53 dummy_5 IN_M 2.82f
C54 m11m12 bias21 0.836f
C55 m3m4 dummy_3 2.84f
C56 VCC m1_44990_37960# 31.6f
C57 VCC IB 27.6f
C58 OUT VB_B 5.56f
C59 m11m12 dummy_3 20.7f
C60 dummy_2 OUT 15.7f
C61 m11m12 m3m4 0.403f
C62 m9m10 m1m2 0.118p
C63 bias21 m1_44990_37960# 1.69f
C64 bias21 IB 0.619f
C65 VCC m1m2 0.153p
C66 IN_P m1_44990_37960# 13.5f
C67 bias3 VB_B 0.977f
C68 bias1 m1m2 61.6f
C69 m9m10 dummy_9 35.8f
C70 dummy_5 bias3 0.399f
C71 IN_M bias3 10.4f
C72 dummy_9 VCC 0.126p
C73 VB_A m1m2 6.26f
C74 VCC VB_B 4.16f
C75 dummy_2 m9m10 2.69f
C76 dummy_2 VCC 13f
C77 VCC dummy_5 11.7f
C78 OUT bias3 0.977f
C79 bias1 dummy_9 0.106p
C80 VCC IN_M 12.8f
C81 bias1 VB_B 5.61f
C82 dummy_4 VSS 3.54f
C83 bias21 VSS 17.4f
C84 OUT VSS 27.3f
C85 m11m12 VSS 24.7f
C86 dummy_5 VSS 17.1f
C87 IN_P VSS 13.3f
C88 VCC VSS 22.5p
C89 dummy_9 VSS 0.175p
C90 bias1 VSS 3.62p
C91 m9m10 VSS 0.169p
C92 dummy_2 VSS 25.9f
C93 VB_A VSS 0.1p
C94 bias3 VSS 45.7f
C95 m1_44990_37960# VSS 9.49f
C96 IN_M VSS 9.08f
C97 m3m4 VSS 19.9f
C98 m1m2 VSS 0.157p
C99 dummy_3 VSS 43.3f
C100 VB_B VSS 0.19p
C101 dummy_100 VSS 8.79f
C102 IB VSS 23.4f
.ends

