magic
tech sky130A
magscale 1 2
timestamp 1697746166
<< nwell >>
rect 60000 90000 106000 144400
rect 38000 16600 106000 90000
rect 38000 16200 65000 16600
rect 65120 16200 65660 16600
rect 65800 16200 106000 16600
rect 38000 14000 106000 16200
<< pwell >>
rect 40000 91600 56800 139000
<< pmos >>
rect 43900 86600 44060 87220
<< psubdiff >>
rect 40300 134600 40460 134660
rect 42120 134600 42380 134660
rect 40300 134460 40460 134520
rect 42120 134460 42380 134520
rect 40300 134340 40460 134400
rect 42120 134340 42380 134400
rect 40300 134200 40460 134260
rect 42120 134200 42380 134260
rect 40300 134040 40460 134100
rect 42120 134040 42380 134100
<< nsubdiff >>
rect 60140 143840 60260 143880
rect 60740 143840 60860 143880
rect 60140 143720 60260 143760
rect 60740 143720 60860 143760
rect 60140 143600 60260 143640
rect 60740 143600 60860 143640
rect 60140 143460 60260 143500
rect 60740 143460 60860 143500
rect 60140 143320 60260 143360
rect 60740 143320 60860 143360
<< psubdiffcont >>
rect 40460 134600 42120 134660
rect 40460 134460 42120 134520
rect 40460 134340 42120 134400
rect 40460 134200 42120 134260
rect 40460 134040 42120 134100
<< nsubdiffcont >>
rect 60260 143840 60740 143880
rect 60260 143720 60740 143760
rect 60260 143600 60740 143640
rect 60260 143460 60740 143500
rect 60260 143320 60740 143360
<< locali >>
rect 40300 134600 40460 134660
rect 42120 134600 42380 134660
rect 40300 134460 40460 134520
rect 42120 134460 42380 134520
rect 40300 134340 40460 134400
rect 42120 134340 42380 134400
rect 40300 134200 40460 134260
rect 42120 134200 42380 134260
rect 40300 134040 40460 134100
rect 42120 134040 42380 134100
<< viali >>
rect 60140 143840 60260 143880
rect 60260 143840 60740 143880
rect 60740 143840 60860 143880
rect 60140 143760 60860 143840
rect 60140 143720 60260 143760
rect 60260 143720 60740 143760
rect 60740 143720 60860 143760
rect 60140 143640 60860 143720
rect 60140 143600 60260 143640
rect 60260 143600 60740 143640
rect 60740 143600 60860 143640
rect 60140 143500 60860 143600
rect 60140 143460 60260 143500
rect 60260 143460 60740 143500
rect 60740 143460 60860 143500
rect 60140 143360 60860 143460
rect 60140 143320 60260 143360
rect 60260 143320 60740 143360
rect 60740 143320 60860 143360
rect 40460 134600 42120 134660
rect 40460 134520 42120 134600
rect 40460 134460 42120 134520
rect 40460 134400 42120 134460
rect 40460 134340 42120 134400
rect 40460 134260 42120 134340
rect 40460 134200 42120 134260
rect 40460 134100 42120 134200
rect 40460 134040 42120 134100
<< metal1 >>
rect 58190 143400 58200 144400
rect 59200 143880 68400 144400
rect 59200 143400 60140 143880
rect 60128 143320 60140 143400
rect 60860 143400 68400 143880
rect 69600 143400 75600 144400
rect 76600 143400 82800 144400
rect 84000 143400 90000 144400
rect 91200 143400 97200 144400
rect 60860 143320 60872 143400
rect 60128 143314 60872 143320
rect 62990 142200 63000 143000
rect 64000 142200 64010 143000
rect 66600 142988 67600 143000
rect 61900 141780 62000 141800
rect 40400 134660 42200 134800
rect 40400 134040 40460 134660
rect 42120 134040 42200 134660
rect 40400 133800 42200 134040
rect 40390 133000 40400 133800
rect 42200 133000 42210 133800
rect 42200 131600 51400 132000
rect 41190 129800 41200 130200
rect 41600 129800 41610 130200
rect 41200 37200 41600 129800
rect 42200 37600 42600 131600
rect 48720 131170 48800 131200
rect 48670 131110 48680 131170
rect 48840 131110 48850 131170
rect 49040 131110 49050 131170
rect 49230 131110 49240 131170
rect 49420 131120 49430 131180
rect 49610 131120 49620 131180
rect 49800 131120 49810 131180
rect 49990 131120 50000 131180
rect 50620 131170 50700 131200
rect 50180 131110 50190 131170
rect 50370 131110 50380 131170
rect 50560 131110 50570 131170
rect 50750 131110 50760 131170
rect 48600 131000 48630 131080
rect 48600 130900 48610 131000
rect 48670 130900 48680 131000
rect 48170 130360 48180 130600
rect 48420 130360 48430 130600
rect 48180 116800 48420 130360
rect 48600 128650 48630 130900
rect 48720 130800 48800 131110
rect 48890 131000 48920 131080
rect 50500 131000 50530 131090
rect 48830 130900 48840 131000
rect 48900 130900 48920 131000
rect 48980 130900 48990 131000
rect 49050 130900 49060 131000
rect 49200 130900 49210 131000
rect 49280 130900 49290 131000
rect 49360 130900 49370 131000
rect 49440 130900 49450 131000
rect 49580 130900 49590 131000
rect 49660 130900 49670 131000
rect 49740 130900 49750 131000
rect 49820 130900 49830 131000
rect 49960 130900 49970 131000
rect 50040 130900 50050 131000
rect 50130 130900 50140 131000
rect 50210 130900 50220 131000
rect 50340 130900 50350 131000
rect 50420 130900 50430 131000
rect 50500 130900 50510 131000
rect 50580 130900 50590 131000
rect 48660 130740 48670 130800
rect 48850 130740 48860 130800
rect 48720 128830 48800 130740
rect 48660 128770 48670 128830
rect 48850 128770 48860 128830
rect 48720 128740 48800 128770
rect 48590 128550 48600 128650
rect 48670 128550 48680 128650
rect 48600 128490 48630 128550
rect 48720 128510 48790 128740
rect 48890 128660 48920 130900
rect 49040 130740 49050 130800
rect 49230 130740 49240 130800
rect 49420 130750 49430 130810
rect 49610 130750 49620 130810
rect 49800 130750 49810 130810
rect 49990 130750 50000 130810
rect 50180 130740 50190 130800
rect 50370 130740 50380 130800
rect 48960 130360 48970 130460
rect 49070 130360 49080 130460
rect 48970 129920 49010 130360
rect 49270 130300 49310 130310
rect 49240 130240 49250 130300
rect 49310 130240 49320 130300
rect 49040 130000 49050 130070
rect 49220 130000 49230 130070
rect 49120 128920 49150 129990
rect 49270 129920 49310 130240
rect 49350 128920 49390 130630
rect 49500 128920 49540 130690
rect 49650 130300 49760 130630
rect 49650 130230 49670 130300
rect 49740 130230 49760 130300
rect 49650 128950 49760 130230
rect 49880 128920 49920 130690
rect 50030 130050 50070 130630
rect 50340 130370 50350 130470
rect 50450 130370 50460 130470
rect 50010 130000 50070 130050
rect 50030 128920 50070 130000
rect 50100 130300 50140 130310
rect 50100 130240 50110 130300
rect 50170 130240 50180 130300
rect 50100 129920 50140 130240
rect 50180 130000 50190 130070
rect 50360 130000 50370 130070
rect 50260 128920 50290 129990
rect 50410 129920 50450 130370
rect 49040 128890 49620 128920
rect 49800 128890 50380 128920
rect 49040 128770 49050 128830
rect 49230 128770 49240 128830
rect 49420 128770 49430 128830
rect 49610 128770 49620 128830
rect 49800 128770 49810 128830
rect 49990 128770 50000 128830
rect 50180 128770 50190 128830
rect 50370 128770 50380 128830
rect 50500 128660 50530 130900
rect 50620 130800 50700 131110
rect 50790 131000 50820 131080
rect 50730 130900 50740 131000
rect 50810 130900 50820 131000
rect 50560 130740 50570 130800
rect 50750 130740 50760 130800
rect 50620 128830 50700 130740
rect 50560 128770 50570 128830
rect 50750 128770 50760 128830
rect 50620 128740 50700 128770
rect 48820 128560 48830 128660
rect 48900 128560 48920 128660
rect 48990 128560 49000 128660
rect 49070 128560 49080 128660
rect 49200 128560 49210 128660
rect 49280 128560 49290 128660
rect 49370 128560 49380 128660
rect 49450 128560 49460 128660
rect 49580 128560 49590 128660
rect 49660 128560 49670 128660
rect 49750 128560 49760 128660
rect 49830 128560 49840 128660
rect 49960 128560 49970 128660
rect 50040 128560 50050 128660
rect 50130 128560 50140 128660
rect 50210 128560 50220 128660
rect 50340 128560 50350 128660
rect 50420 128560 50430 128660
rect 50500 128560 50520 128660
rect 50590 128560 50600 128660
rect 48720 128460 48800 128510
rect 48890 128490 48920 128560
rect 50500 128500 50530 128560
rect 50630 128490 50690 128740
rect 50790 128660 50820 130900
rect 51200 130200 51400 131600
rect 51710 130360 51720 130600
rect 51960 130360 51970 130600
rect 51190 130000 51200 130200
rect 51400 130000 51410 130200
rect 50720 128560 50730 128660
rect 50800 128560 50820 128660
rect 50790 128490 50820 128560
rect 50620 128460 50700 128490
rect 48660 128400 48670 128460
rect 48850 128400 48860 128460
rect 49040 128400 49050 128460
rect 49230 128400 49240 128460
rect 49420 128400 49430 128460
rect 49610 128400 49620 128460
rect 49800 128400 49810 128460
rect 49990 128400 50000 128460
rect 50180 128400 50190 128460
rect 50370 128400 50380 128460
rect 50560 128400 50570 128460
rect 50750 128400 50760 128460
rect 48180 116640 48200 116800
rect 48190 116600 48200 116640
rect 48400 116640 48420 116800
rect 48400 116600 48410 116640
rect 51720 114880 51960 130360
rect 44880 114780 51960 114880
rect 43790 112900 43800 113300
rect 44400 112900 44410 113300
rect 43490 112360 43630 112660
rect 43490 111860 43620 112360
rect 43720 111860 43730 112360
rect 43490 92820 43630 111860
rect 43490 92320 43620 92820
rect 43720 92320 43730 92820
rect 43490 92080 43630 92320
rect 43800 92000 44400 112900
rect 44590 111860 44600 112360
rect 44700 111860 44710 112360
rect 44760 111620 44840 112440
rect 44880 112402 44960 114780
rect 48190 113900 48200 114000
rect 46280 113820 48200 113900
rect 45290 112900 45300 113300
rect 45900 112900 45910 113300
rect 44880 111704 44962 112402
rect 45010 111860 45020 112360
rect 45120 111860 45130 112360
rect 44880 111620 44960 111704
rect 44756 111516 44830 111620
rect 44690 92820 44830 111516
rect 44890 111526 44960 111620
rect 44890 93280 45030 111526
rect 44880 92896 44960 93280
rect 44590 92320 44600 92820
rect 44700 92320 44830 92820
rect 45010 92340 45020 92840
rect 45120 92340 45130 92840
rect 44690 92080 44830 92320
rect 45300 92000 45900 112900
rect 45990 111860 46000 112360
rect 46100 111860 46110 112360
rect 46160 111620 46240 112380
rect 46280 111620 46360 113820
rect 48190 113800 48200 113820
rect 48400 113900 48410 114000
rect 48400 113820 49040 113900
rect 48400 113800 48410 113820
rect 46690 112900 46700 113300
rect 47300 112900 47310 113300
rect 48090 112900 48100 113300
rect 48700 112900 48710 113300
rect 46410 111860 46420 112360
rect 46520 111860 46530 112360
rect 46160 111526 46230 111620
rect 46090 93280 46230 111526
rect 46290 111532 46362 111620
rect 46290 93280 46430 111532
rect 45990 92340 46000 92840
rect 46100 92340 46110 92840
rect 46160 91200 46240 93280
rect 46280 92080 46360 93280
rect 46410 92340 46420 92840
rect 46520 92340 46530 92840
rect 46700 92000 47300 112900
rect 47390 111860 47400 112360
rect 47500 111860 47510 112360
rect 47560 111638 47760 112380
rect 47810 111860 47820 112360
rect 47920 111860 47930 112360
rect 47570 111620 47760 111638
rect 47570 111536 47762 111620
rect 47570 111534 47830 111536
rect 47490 93280 47830 111534
rect 47390 92340 47400 92840
rect 47500 92340 47510 92840
rect 47560 91760 47760 93280
rect 47810 92340 47820 92840
rect 47940 92340 47950 92840
rect 48100 92000 48700 112900
rect 48790 111860 48800 112360
rect 48900 111860 48910 112360
rect 48960 111624 49040 113820
rect 49490 112900 49500 113300
rect 50100 112900 50110 113300
rect 48962 111620 49040 111624
rect 49080 111620 49160 112360
rect 49210 111860 49220 112360
rect 49320 111860 49330 112360
rect 48962 111514 49030 111620
rect 48890 93300 49030 111514
rect 49090 111512 49162 111620
rect 49090 93300 49230 111512
rect 48890 93280 49040 93300
rect 48790 92340 48800 92840
rect 48900 92340 48910 92840
rect 48960 92100 49040 93280
rect 49080 93280 49230 93300
rect 47550 91460 47560 91760
rect 47760 91460 47770 91760
rect 46000 90800 46400 91200
rect 49080 91000 49160 93280
rect 49210 92340 49220 92840
rect 49320 92340 49330 92840
rect 49500 92000 50100 112900
rect 50360 112360 50432 114780
rect 50480 114766 50560 114780
rect 50890 112900 50900 113300
rect 51500 112900 51510 113300
rect 50190 111860 50200 112360
rect 50300 111860 50310 112360
rect 50360 111628 50440 112360
rect 50366 111620 50440 111628
rect 50480 111632 50560 112314
rect 50610 111860 50620 112360
rect 50720 111860 50730 112360
rect 50480 111620 50558 111632
rect 50366 111518 50430 111620
rect 50290 93300 50430 111518
rect 50490 111522 50558 111620
rect 50490 93300 50630 111522
rect 50290 93280 50440 93300
rect 50190 92340 50200 92840
rect 50300 92340 50310 92840
rect 50360 92100 50440 93280
rect 50480 93280 50630 93300
rect 50480 92766 50560 93280
rect 50610 92766 50620 92840
rect 50720 92766 50730 92840
rect 50480 92388 50516 92766
rect 50726 92388 50736 92766
rect 50480 92100 50560 92388
rect 50610 92340 50620 92388
rect 50720 92340 50730 92388
rect 50900 92000 51500 112900
rect 51690 112360 51830 112660
rect 51590 111860 51600 112360
rect 51700 111860 51830 112360
rect 51690 92840 51830 111860
rect 51590 92340 51600 92840
rect 51700 92340 51830 92840
rect 51690 92070 51830 92340
rect 45990 90400 46000 90800
rect 46400 90400 46410 90800
rect 46000 88760 46400 90400
rect 49000 88760 49200 91000
rect 44920 88540 50460 88760
rect 43890 87500 43900 87900
rect 44500 87500 44510 87900
rect 43580 66480 43660 87300
rect 43820 86660 43830 87040
rect 43820 66820 43830 67220
rect 43900 66400 44500 87500
rect 44570 86660 44580 87040
rect 44610 66820 44620 67200
rect 44720 66480 44800 87300
rect 44920 86060 44980 88540
rect 46320 88020 47560 88340
rect 47760 88020 49060 88340
rect 45290 87500 45300 87900
rect 45900 87500 45910 87900
rect 45050 86660 45060 87040
rect 45160 86660 45170 87040
rect 44920 67720 45060 86060
rect 44920 66180 44980 67720
rect 45050 66820 45060 67200
rect 45220 66820 45230 67200
rect 45300 66400 45900 87500
rect 46030 86660 46040 87040
rect 46140 86660 46150 87040
rect 46200 86080 46260 87320
rect 46120 67720 46260 86080
rect 45950 66820 45960 67200
rect 46120 66820 46130 67200
rect 46200 66540 46260 67720
rect 46320 86060 46380 88020
rect 46690 87500 46700 87900
rect 47300 87500 47310 87900
rect 48090 87500 48100 87900
rect 48700 87500 48710 87900
rect 46450 86660 46460 87040
rect 46620 86660 46630 87040
rect 46320 67720 46460 86060
rect 46190 66440 46200 66540
rect 46260 66440 46270 66540
rect 46200 66420 46260 66440
rect 46320 66420 46380 67720
rect 46450 66820 46460 67200
rect 46600 66820 46610 67200
rect 46700 66400 47300 87500
rect 47410 86660 47420 87040
rect 47520 86660 47530 87040
rect 47600 86060 47780 87380
rect 47850 86660 47860 87060
rect 48020 86660 48030 87060
rect 47520 67720 47860 86060
rect 47370 66820 47380 67200
rect 47520 66820 47530 67200
rect 47600 66200 47780 67720
rect 47850 66820 47860 67200
rect 48000 66820 48010 67200
rect 48100 66400 48700 87500
rect 48810 86660 48820 87040
rect 48940 86660 48950 87040
rect 49000 86060 49060 88020
rect 49490 87500 49500 87900
rect 50100 87500 50110 87900
rect 48920 67720 49060 86060
rect 48810 66820 48820 67200
rect 48940 66820 48950 67200
rect 49000 66440 49060 67720
rect 49120 86060 49180 87300
rect 49250 86660 49260 87040
rect 49420 86660 49430 87040
rect 49120 67720 49260 86060
rect 49120 66540 49180 67720
rect 49250 66820 49260 67200
rect 49380 66820 49390 67200
rect 49110 66440 49120 66540
rect 49180 66440 49190 66540
rect 49500 66400 50100 87500
rect 50170 86660 50180 87040
rect 50320 86660 50330 87040
rect 50400 86060 50460 88540
rect 50890 87500 50900 87900
rect 51500 87500 51510 87900
rect 50320 67720 50460 86060
rect 50210 66820 50220 67200
rect 50340 66820 50350 67200
rect 50400 66460 50460 67720
rect 50580 66460 50660 87300
rect 50800 86660 50810 87040
rect 50760 66820 50770 67200
rect 50900 66400 51500 87500
rect 51720 87040 51800 87300
rect 51590 86660 51600 87040
rect 51740 86660 51800 87040
rect 51610 66820 51620 67200
rect 51720 66480 51800 86660
rect 47600 65800 60500 66200
rect 46020 54640 50760 54680
rect 44990 51800 45000 52200
rect 45400 51800 45410 52200
rect 45000 38480 45400 51800
rect 46020 47820 46060 54640
rect 46190 54300 46200 54500
rect 46600 54300 46610 54500
rect 46200 47900 46600 54300
rect 46740 54060 46860 54640
rect 46990 54300 47000 54500
rect 47400 54300 47410 54500
rect 46740 54040 46880 54060
rect 46720 53060 46880 54040
rect 46720 49100 46760 53060
rect 46820 52800 46860 52840
rect 46810 51820 46820 52800
rect 46920 51820 46930 52800
rect 46820 49220 46860 51820
rect 46720 47820 46860 49100
rect 47000 47900 47400 54300
rect 47520 53060 47660 54640
rect 47790 54300 47800 54500
rect 48200 54300 48210 54500
rect 47520 51620 47560 52840
rect 47620 51800 47660 53060
rect 47520 50340 47660 51620
rect 47510 49320 47520 50340
rect 47660 49320 47670 50340
rect 47520 49220 47660 49320
rect 47520 47820 47660 49120
rect 47800 47900 48200 54300
rect 48320 51800 48460 54640
rect 48590 54300 48600 54500
rect 49000 54300 49010 54500
rect 48320 51580 48460 51620
rect 48310 50560 48320 51580
rect 48460 50560 48470 51580
rect 48320 49220 48460 50560
rect 48320 47820 48460 49120
rect 48600 47900 49000 54300
rect 49120 53060 49260 54640
rect 49390 54300 49400 54500
rect 49800 54300 49810 54500
rect 49120 51800 49160 53060
rect 49120 50340 49160 51620
rect 49220 50340 49260 52840
rect 49110 49320 49120 50340
rect 49260 49320 49270 50340
rect 49120 49220 49160 49320
rect 49220 49220 49260 49320
rect 49120 47820 49260 49120
rect 49400 47900 49800 54300
rect 49920 53060 50060 54640
rect 50190 54300 50200 54500
rect 50600 54300 50610 54500
rect 49920 52800 49960 52860
rect 49850 51820 49860 52800
rect 49960 51820 49970 52800
rect 49920 49240 49960 51820
rect 50020 49240 50060 53060
rect 49920 47820 50060 49120
rect 50200 47900 50600 54300
rect 50720 47820 50760 54640
rect 46020 47780 50760 47820
rect 44990 37960 45000 38480
rect 45400 37960 45410 38480
rect 42200 37400 51300 37600
rect 51520 37400 51600 37600
rect 41200 37000 50100 37200
rect 50320 37000 50400 37200
rect 49040 36720 52580 36780
rect 49040 35640 49140 36720
rect 49190 35700 49200 35800
rect 49400 35700 52200 35800
rect 52400 35700 52410 35800
rect 52480 35640 52580 36720
rect 49040 35580 52580 35640
rect 49040 35480 49380 35580
rect 49870 35480 49880 35540
rect 49940 35480 49950 35540
rect 50470 35480 50480 35540
rect 50540 35480 50550 35540
rect 51070 35480 51080 35540
rect 51140 35480 51150 35540
rect 51670 35480 51680 35540
rect 51740 35480 51750 35540
rect 52240 35480 52580 35580
rect 49040 34400 49140 35480
rect 49490 35240 49500 35380
rect 49720 35240 49730 35380
rect 50090 35240 50100 35380
rect 50320 35240 50330 35380
rect 50690 35240 50700 35380
rect 50920 35240 50930 35380
rect 51290 35240 51300 35380
rect 51520 35240 51530 35380
rect 51890 35240 51900 35380
rect 52120 35240 52130 35380
rect 49500 34600 49724 35240
rect 50100 34600 50320 35240
rect 50700 34600 50924 35240
rect 51300 34600 51524 35240
rect 51900 34600 52124 35240
rect 49190 34500 49200 34600
rect 49400 34500 49410 34600
rect 49500 34500 49860 34600
rect 49960 34500 50460 34600
rect 50560 34500 51060 34600
rect 51160 34500 51660 34600
rect 51760 34500 52124 34600
rect 52190 34500 52200 34600
rect 52400 34500 52410 34600
rect 49040 34240 49380 34400
rect 49040 33160 49140 34240
rect 49500 33400 49724 34500
rect 49870 34240 49880 34400
rect 49940 34240 49950 34400
rect 50100 33400 50320 34500
rect 50470 34240 50480 34400
rect 50540 34240 50550 34400
rect 50700 33400 50924 34500
rect 51070 34240 51080 34400
rect 51140 34240 51150 34400
rect 51300 33400 51524 34500
rect 51670 34240 51680 34400
rect 51740 34240 51750 34400
rect 51900 33400 52124 34500
rect 52480 34400 52580 35480
rect 52240 34240 52580 34400
rect 49190 33300 49200 33400
rect 49400 33300 49410 33400
rect 49500 33300 49880 33400
rect 49960 33300 50460 33400
rect 50560 33300 51060 33400
rect 51160 33300 51660 33400
rect 51760 33300 52124 33400
rect 52190 33300 52200 33400
rect 52400 33300 52410 33400
rect 49040 33020 49380 33160
rect 49040 31940 49140 33020
rect 49500 32100 49724 33300
rect 49870 33000 49880 33160
rect 49940 33000 49950 33160
rect 50100 32100 50320 33300
rect 50470 33000 50480 33160
rect 50540 33000 50550 33160
rect 50700 32100 50924 33300
rect 51070 33000 51080 33160
rect 51140 33000 51150 33160
rect 51300 32100 51524 33300
rect 51670 33000 51680 33160
rect 51740 33000 51750 33160
rect 51900 32100 52124 33300
rect 52480 33160 52580 34240
rect 52240 33020 52580 33160
rect 49190 32000 49200 32100
rect 49400 32000 49410 32100
rect 49500 32000 49860 32100
rect 49960 32000 50460 32100
rect 50560 32000 51060 32100
rect 51160 32000 51660 32100
rect 51760 32000 52124 32100
rect 52190 32000 52200 32100
rect 52400 32000 52410 32100
rect 49040 31780 49380 31940
rect 49040 30700 49140 31780
rect 49500 30900 49724 32000
rect 49870 31780 49880 31940
rect 49940 31780 49950 31940
rect 50100 30900 50320 32000
rect 50470 31780 50480 31940
rect 50540 31780 50550 31940
rect 50700 30900 50924 32000
rect 51070 31780 51080 31940
rect 51140 31780 51150 31940
rect 51300 30900 51524 32000
rect 51670 31780 51680 31940
rect 51740 31780 51750 31940
rect 51900 30900 52124 32000
rect 52480 31940 52580 33020
rect 52240 31780 52580 31940
rect 49190 30800 49200 30900
rect 49400 30800 49410 30900
rect 49500 30800 49880 30900
rect 49960 30800 50460 30900
rect 50560 30800 51060 30900
rect 51160 30800 51660 30900
rect 51760 30800 52124 30900
rect 52190 30800 52200 30900
rect 52400 30800 52410 30900
rect 49040 30540 49380 30700
rect 49040 29460 49140 30540
rect 49500 29700 49724 30800
rect 49870 30540 49880 30700
rect 49940 30540 49950 30700
rect 50100 29700 50320 30800
rect 50470 30540 50480 30700
rect 50540 30540 50550 30700
rect 50700 29700 50924 30800
rect 51070 30540 51080 30700
rect 51140 30540 51150 30700
rect 51300 29700 51524 30800
rect 51670 30540 51680 30700
rect 51740 30540 51750 30700
rect 51900 29700 52124 30800
rect 52480 30700 52580 31780
rect 52240 30540 52580 30700
rect 49190 29600 49200 29700
rect 49400 29600 49410 29700
rect 49500 29600 49880 29700
rect 49960 29600 50460 29700
rect 50560 29600 51060 29700
rect 51160 29600 51660 29700
rect 51760 29600 52124 29700
rect 52190 29600 52200 29700
rect 52400 29600 52410 29700
rect 49040 29300 49380 29460
rect 49040 28220 49140 29300
rect 49500 28500 49724 29600
rect 49870 29300 49880 29460
rect 49940 29300 49950 29460
rect 50100 28500 50320 29600
rect 50470 29300 50480 29460
rect 50540 29300 50550 29460
rect 50700 28500 50924 29600
rect 51070 29300 51080 29460
rect 51140 29300 51150 29460
rect 51300 28500 51524 29600
rect 51670 29300 51680 29460
rect 51740 29300 51750 29460
rect 51900 28500 52124 29600
rect 52480 29460 52580 30540
rect 52240 29300 52580 29460
rect 49190 28400 49200 28500
rect 49400 28400 49410 28500
rect 49500 28400 49880 28500
rect 49960 28400 50460 28500
rect 50560 28400 51060 28500
rect 51160 28400 51660 28500
rect 51760 28400 52124 28500
rect 52190 28400 52200 28500
rect 52400 28400 52410 28500
rect 49040 28060 49380 28220
rect 49040 26980 49140 28060
rect 49500 27200 49724 28400
rect 49870 28080 49880 28220
rect 49940 28080 49950 28220
rect 50100 27200 50320 28400
rect 50470 28080 50480 28220
rect 50540 28080 50550 28220
rect 50700 27200 50924 28400
rect 51070 28080 51080 28220
rect 51140 28080 51150 28220
rect 51300 27200 51524 28400
rect 51670 28080 51680 28220
rect 51740 28080 51750 28220
rect 51900 27200 52124 28400
rect 52480 28220 52580 29300
rect 52240 28060 52580 28220
rect 49190 27100 49200 27200
rect 49400 27100 49410 27200
rect 49500 27100 49880 27200
rect 49960 27100 50460 27200
rect 50560 27100 51060 27200
rect 51160 27100 51660 27200
rect 51760 27100 52124 27200
rect 52190 27100 52200 27200
rect 52400 27100 52410 27200
rect 49040 26820 49380 26980
rect 49040 25760 49140 26820
rect 49500 26000 49724 27100
rect 49870 26820 49880 26980
rect 49940 26820 49950 26980
rect 50100 26000 50320 27100
rect 50470 26840 50480 27000
rect 50540 26840 50550 27000
rect 50700 26000 50924 27100
rect 51070 26840 51080 27000
rect 51140 26840 51150 27000
rect 51300 26000 51524 27100
rect 51670 26840 51680 27000
rect 51740 26840 51750 27000
rect 51900 26000 52124 27100
rect 52480 26980 52580 28060
rect 52240 26820 52580 26980
rect 49190 25900 49200 26000
rect 49400 25900 49410 26000
rect 49500 25900 49880 26000
rect 49960 25900 50460 26000
rect 50560 25900 51060 26000
rect 51160 25900 51660 26000
rect 51760 25900 52124 26000
rect 52190 25900 52200 26000
rect 52400 25900 52410 26000
rect 49040 25600 49380 25760
rect 49040 24520 49140 25600
rect 49500 24800 49724 25900
rect 49870 25600 49880 25760
rect 49940 25600 49950 25760
rect 50100 24800 50320 25900
rect 50470 25600 50480 25760
rect 50540 25600 50550 25760
rect 50700 24800 50924 25900
rect 51070 25600 51080 25760
rect 51140 25600 51150 25760
rect 51300 24800 51524 25900
rect 51670 25600 51680 25760
rect 51740 25600 51750 25760
rect 51900 24800 52124 25900
rect 52480 25760 52580 26820
rect 52240 25600 52580 25760
rect 49190 24700 49200 24800
rect 49400 24700 49410 24800
rect 49500 24700 49880 24800
rect 49960 24700 50460 24800
rect 50560 24700 51060 24800
rect 51160 24700 51660 24800
rect 51760 24700 52124 24800
rect 52190 24700 52200 24800
rect 52400 24700 52410 24800
rect 49040 24360 49380 24520
rect 49040 23280 49140 24360
rect 49500 23500 49724 24700
rect 49870 24360 49880 24520
rect 49940 24360 49950 24520
rect 50100 23500 50320 24700
rect 50470 24360 50480 24520
rect 50540 24360 50550 24520
rect 50700 23500 50924 24700
rect 51070 24360 51080 24520
rect 51140 24360 51150 24520
rect 51300 23500 51524 24700
rect 51670 24360 51680 24520
rect 51740 24360 51750 24520
rect 51900 23500 52124 24700
rect 52480 24520 52580 25600
rect 52240 24360 52580 24520
rect 49190 23400 49200 23500
rect 49400 23400 49410 23500
rect 49500 23400 49880 23500
rect 49960 23400 50460 23500
rect 50560 23400 51060 23500
rect 51160 23400 51660 23500
rect 51760 23400 52124 23500
rect 52190 23400 52200 23500
rect 52400 23400 52410 23500
rect 49040 23120 49380 23280
rect 49040 22040 49140 23120
rect 49500 22300 49724 23400
rect 49870 23120 49880 23280
rect 49940 23120 49950 23280
rect 50100 22300 50320 23400
rect 50470 23120 50480 23280
rect 50540 23120 50550 23280
rect 50700 22320 50924 23400
rect 51070 23120 51080 23280
rect 51140 23120 51150 23280
rect 51300 22320 51524 23400
rect 51670 23120 51680 23280
rect 51740 23120 51750 23280
rect 49190 22200 49200 22300
rect 49400 22200 49410 22300
rect 49500 22200 49880 22300
rect 49960 22200 50460 22300
rect 50560 22220 51060 22320
rect 51160 22220 51660 22320
rect 51900 22300 52124 23400
rect 52480 23280 52580 24360
rect 52240 23120 52580 23280
rect 49040 21880 49380 22040
rect 49040 20800 49140 21880
rect 49500 21000 49724 22200
rect 49870 21880 49880 22040
rect 49940 21880 49950 22040
rect 50100 21000 50320 22200
rect 50470 21880 50480 22040
rect 50540 21880 50550 22040
rect 50700 21000 50924 22220
rect 51070 21880 51080 22040
rect 51140 21880 51150 22040
rect 51300 21000 51524 22220
rect 51760 22200 52124 22300
rect 52190 22200 52200 22300
rect 52400 22200 52410 22300
rect 51670 21880 51680 22040
rect 51740 21880 51750 22040
rect 51900 21000 52124 22200
rect 52480 22040 52580 23120
rect 52240 21880 52580 22040
rect 49190 20900 49200 21000
rect 49400 20900 49410 21000
rect 49500 20900 49860 21000
rect 49960 20900 50460 21000
rect 50560 20900 51060 21000
rect 51160 20900 51660 21000
rect 51760 20900 52124 21000
rect 52190 20900 52200 21000
rect 52400 20900 52410 21000
rect 49040 20660 49380 20800
rect 49040 19580 49140 20660
rect 49500 19800 49724 20900
rect 49870 20660 49880 20820
rect 49940 20660 49950 20820
rect 50100 19800 50320 20900
rect 50470 20660 50480 20820
rect 50540 20660 50550 20820
rect 50700 19800 50924 20900
rect 51070 20660 51080 20820
rect 51140 20660 51150 20820
rect 51300 19800 51524 20900
rect 51670 20660 51680 20820
rect 51740 20660 51750 20820
rect 51900 19800 52124 20900
rect 52240 20800 52400 20810
rect 52480 20800 52580 21880
rect 52240 20660 52580 20800
rect 49190 19700 49200 19800
rect 49400 19700 49410 19800
rect 49500 19700 49860 19800
rect 49960 19700 50480 19800
rect 50560 19700 51080 19800
rect 51160 19700 51680 19800
rect 51760 19700 52124 19800
rect 52190 19700 52200 19800
rect 52400 19700 52410 19800
rect 49040 19420 49380 19580
rect 49040 18340 49140 19420
rect 49500 18600 49724 19700
rect 49870 19420 49880 19580
rect 49940 19420 49950 19580
rect 50100 18600 50320 19700
rect 50470 19420 50480 19580
rect 50540 19420 50550 19580
rect 50700 18600 50924 19700
rect 51070 19420 51080 19580
rect 51140 19420 51150 19580
rect 51300 18600 51524 19700
rect 51670 19420 51680 19580
rect 51740 19420 51750 19580
rect 51900 18600 52124 19700
rect 52480 19580 52580 20660
rect 52240 19420 52580 19580
rect 49190 18500 49200 18600
rect 49400 18500 49410 18600
rect 49500 18500 49880 18600
rect 49960 18500 50480 18600
rect 50560 18500 51080 18600
rect 51160 18500 51680 18600
rect 51760 18500 52124 18600
rect 52190 18500 52200 18600
rect 52400 18500 52410 18600
rect 49040 18180 49380 18340
rect 49040 17100 49140 18180
rect 49500 17300 49724 18500
rect 49870 18180 49880 18340
rect 49940 18180 49950 18340
rect 50100 17300 50320 18500
rect 50470 18180 50480 18340
rect 50540 18180 50550 18340
rect 50700 17300 50924 18500
rect 51070 18180 51080 18340
rect 51140 18180 51150 18340
rect 51300 17300 51524 18500
rect 51670 18180 51680 18340
rect 51740 18180 51750 18340
rect 51900 17300 52124 18500
rect 52480 18340 52580 19420
rect 52240 18180 52580 18340
rect 49190 17200 49200 17300
rect 49400 17200 49410 17300
rect 49500 17200 49860 17300
rect 49960 17200 50460 17300
rect 50560 17200 51060 17300
rect 51160 17200 51660 17300
rect 51760 17200 52124 17300
rect 52190 17200 52200 17300
rect 52400 17200 52410 17300
rect 52480 17100 52580 18180
rect 49040 17000 49380 17100
rect 49870 17040 49880 17100
rect 49940 17040 49950 17100
rect 50470 17040 50480 17100
rect 50540 17040 50550 17100
rect 51070 17040 51080 17100
rect 51140 17040 51150 17100
rect 51670 17040 51680 17100
rect 51740 17040 51750 17100
rect 52240 17000 52580 17100
rect 49040 16940 52580 17000
rect 49040 15860 49140 16940
rect 49190 15900 49200 16000
rect 49400 15900 52200 16000
rect 52400 15900 52410 16000
rect 52480 15860 52580 16940
rect 49040 15800 51080 15860
rect 51140 15800 52580 15860
rect 60100 15100 60500 65800
rect 61900 15880 62060 141780
rect 62260 141200 62270 141400
rect 62260 16400 62270 16600
rect 63000 15760 64000 142200
rect 66582 142194 66592 142988
rect 67612 142194 67622 142988
rect 68400 142200 69600 143400
rect 69990 142200 70000 143000
rect 71000 142200 71010 143000
rect 73990 142200 74000 143000
rect 75000 142200 75010 143000
rect 75600 142200 76600 143400
rect 76990 142200 77000 143000
rect 78000 142200 78010 143000
rect 80990 142200 81000 143000
rect 82000 142200 82010 143000
rect 82800 142200 84000 143400
rect 84990 142200 85000 143000
rect 86000 142200 86010 143000
rect 87990 142200 88000 143000
rect 89000 142200 89010 143000
rect 90000 142200 91200 143400
rect 91990 142200 92000 143000
rect 93000 142200 93010 143000
rect 94990 142200 95000 143000
rect 96000 142200 96010 143000
rect 97200 142200 98400 143400
rect 98990 142200 99000 143000
rect 100000 142200 100010 143000
rect 101990 142200 102000 143000
rect 103000 142200 103010 143000
rect 64910 141200 64920 141400
rect 65120 40200 65300 141800
rect 65000 39800 65300 40200
rect 65120 39000 65300 39800
rect 65000 38600 65300 39000
rect 65120 37800 65300 38600
rect 65000 37400 65300 37800
rect 65120 36600 65300 37400
rect 65000 36200 65300 36600
rect 65120 35200 65300 36200
rect 65000 34800 65300 35200
rect 65120 33800 65300 34800
rect 65000 33400 65300 33800
rect 65120 32600 65300 33400
rect 65000 32200 65300 32600
rect 65120 31400 65300 32200
rect 65000 31000 65300 31400
rect 65120 30200 65300 31000
rect 65000 29800 65300 30200
rect 65120 29000 65300 29800
rect 65000 28600 65300 29000
rect 65120 27800 65300 28600
rect 65000 27400 65300 27800
rect 65120 26400 65300 27400
rect 65000 26000 65300 26400
rect 65120 25400 65300 26000
rect 65000 25000 65300 25400
rect 65120 24000 65300 25000
rect 65000 23600 65300 24000
rect 65120 22800 65300 23600
rect 65000 22400 65300 22800
rect 65120 21600 65300 22400
rect 65000 21200 65300 21600
rect 65120 20400 65300 21200
rect 65000 20000 65300 20400
rect 65120 19000 65300 20000
rect 65000 18600 65300 19000
rect 65120 17800 65300 18600
rect 65000 17400 65300 17800
rect 65120 17120 65300 17400
rect 64910 16400 64920 16600
rect 65120 16400 65130 16600
rect 65180 15880 65300 17120
rect 65500 140520 65600 141800
rect 65650 141200 65660 141400
rect 65860 141200 65870 141400
rect 65500 40200 65660 140520
rect 65500 39800 65800 40200
rect 65500 39000 65660 39800
rect 65500 38600 65800 39000
rect 65500 37800 65660 38600
rect 65500 37400 65800 37800
rect 65500 36600 65660 37400
rect 65500 36200 65800 36600
rect 65500 35200 65660 36200
rect 65500 34800 65800 35200
rect 65500 33800 65660 34800
rect 65500 33400 65800 33800
rect 65500 32600 65660 33400
rect 65500 32200 65800 32600
rect 65500 31400 65660 32200
rect 65500 31000 65800 31400
rect 65500 30200 65660 31000
rect 65500 29800 65800 30200
rect 65500 29000 65660 29800
rect 65500 28600 65800 29000
rect 65500 27800 65660 28600
rect 65500 27400 65800 27800
rect 65500 26400 65660 27400
rect 65500 26000 65800 26400
rect 65500 25400 65660 26000
rect 65500 25000 65800 25400
rect 65500 24000 65660 25000
rect 65500 23600 65800 24000
rect 65500 22800 65660 23600
rect 65500 22400 65800 22800
rect 65500 21600 65660 22400
rect 65500 21200 65800 21600
rect 65500 20400 65660 21200
rect 65500 20000 65800 20400
rect 65500 19000 65660 20000
rect 65500 18600 65800 19000
rect 65500 17800 65660 18600
rect 65500 17400 65800 17800
rect 65500 17120 65660 17400
rect 65500 15100 65600 17120
rect 65650 16400 65660 16600
rect 65860 16400 65870 16600
rect 66600 15760 67600 142194
rect 68800 141800 69200 142200
rect 68780 141600 69200 141800
rect 68510 141200 68520 141400
rect 68720 141200 68730 141400
rect 68780 140560 68900 141600
rect 68720 17120 68900 140560
rect 68510 16400 68520 16600
rect 68720 16400 68730 16600
rect 68780 15600 68900 17120
rect 69100 140520 69200 141600
rect 69250 141200 69260 141400
rect 69460 141200 69470 141400
rect 69100 17120 69260 140520
rect 69100 15600 69200 17120
rect 69250 16400 69260 16600
rect 69460 16400 69470 16600
rect 70000 15780 71000 142200
rect 72110 141200 72120 141400
rect 72320 141200 72330 141400
rect 72380 140540 72500 141800
rect 72320 17120 72500 140540
rect 72110 16400 72120 16600
rect 72320 16400 72330 16600
rect 68780 15300 69200 15600
rect 72380 15400 72500 17120
rect 72700 140520 72800 141800
rect 72850 141200 72860 141400
rect 73060 141200 73070 141400
rect 72700 17120 72860 140520
rect 72380 15300 72400 15400
rect 72500 15300 72510 15400
rect 72700 15100 72800 17120
rect 72850 16400 72860 16600
rect 73060 16400 73070 16600
rect 74000 15780 75000 142200
rect 76000 141800 76400 142200
rect 75710 141200 75720 141400
rect 75920 141200 75930 141400
rect 75980 140520 76100 141800
rect 75920 17120 76100 140520
rect 75710 16400 75720 16600
rect 75920 16400 75930 16600
rect 75980 15600 76100 17120
rect 76300 140520 76400 141800
rect 76450 141200 76460 141400
rect 76660 141200 76670 141400
rect 76300 17120 76460 140520
rect 76300 15600 76400 17120
rect 76450 16400 76460 16600
rect 76660 16400 76670 16600
rect 77000 15780 78000 142200
rect 79310 141200 79320 141400
rect 79520 141200 79530 141400
rect 79600 140520 79700 141800
rect 79520 17120 79700 140520
rect 79310 16400 79320 16600
rect 79520 16400 79530 16600
rect 75980 15300 76400 15600
rect 79580 15400 79700 17120
rect 79900 140520 80000 141800
rect 80050 141200 80060 141400
rect 80260 141200 80270 141400
rect 79900 17120 80060 140520
rect 79580 15300 79600 15400
rect 79700 15300 79710 15400
rect 79900 15100 80000 17120
rect 80050 16400 80060 16600
rect 80260 16400 80270 16600
rect 81000 15780 82000 142200
rect 83200 141800 83600 142200
rect 82910 141200 82920 141400
rect 83120 141200 83130 141400
rect 83200 140520 83300 141800
rect 83120 17120 83300 140520
rect 82910 16400 82920 16600
rect 83120 16400 83130 16600
rect 83180 15600 83300 17120
rect 83500 140520 83600 141800
rect 83650 141200 83660 141400
rect 83860 141200 83870 141400
rect 83500 17120 83660 140520
rect 83500 15600 83600 17120
rect 83650 16400 83660 16600
rect 83860 16400 83870 16600
rect 85000 15780 86000 142200
rect 86510 141200 86520 141400
rect 86720 141200 86730 141400
rect 86800 140520 86900 141800
rect 86720 17120 86900 140520
rect 86510 16400 86520 16600
rect 86720 16400 86730 16600
rect 83180 15300 83600 15600
rect 86780 15400 86900 17120
rect 87100 140520 87200 141800
rect 87250 141200 87260 141400
rect 87460 141200 87470 141400
rect 87100 17120 87260 140520
rect 86780 15300 86800 15400
rect 86900 15300 86910 15400
rect 87100 15100 87200 17120
rect 87250 16400 87260 16600
rect 87460 16400 87470 16600
rect 88000 15780 89000 142200
rect 90400 141800 90800 142200
rect 90110 141200 90120 141400
rect 90320 141200 90330 141400
rect 90400 140520 90500 141800
rect 90320 17120 90500 140520
rect 90110 16400 90120 16600
rect 90320 16400 90330 16600
rect 90380 15600 90500 17120
rect 90700 140520 90800 141800
rect 90850 141200 90860 141400
rect 91060 141200 91070 141400
rect 90700 17120 90860 140520
rect 90700 15600 90800 17120
rect 90850 16400 90860 16600
rect 91060 16400 91070 16600
rect 92000 15780 93000 142200
rect 93710 141200 93720 141400
rect 93920 141200 93930 141400
rect 94000 140520 94100 141800
rect 93920 17120 94100 140520
rect 93710 16400 93720 16600
rect 93920 16400 93930 16600
rect 90380 15300 90800 15600
rect 93980 15400 94100 17120
rect 94300 140520 94400 141800
rect 94450 141200 94460 141400
rect 94660 141200 94670 141400
rect 94300 17120 94460 140520
rect 93980 15300 94000 15400
rect 94100 15300 94110 15400
rect 94300 15100 94400 17120
rect 94450 16400 94460 16600
rect 94660 16400 94670 16600
rect 95000 15780 96000 142200
rect 97600 141800 98000 142200
rect 97310 141200 97320 141400
rect 97520 141200 97530 141400
rect 97600 140520 97700 141800
rect 97520 17120 97700 140520
rect 97310 16400 97320 16600
rect 97520 16400 97530 16600
rect 97580 15600 97700 17120
rect 97900 140520 98000 141800
rect 98050 141200 98060 141400
rect 98260 141200 98270 141400
rect 97900 17120 98060 140520
rect 97900 15600 98000 17120
rect 98050 16400 98060 16600
rect 98260 16400 98270 16600
rect 99000 15780 100000 142200
rect 100910 141200 100920 141400
rect 101120 141200 101130 141400
rect 101200 140520 101300 141800
rect 101120 17120 101300 140520
rect 100910 16400 100920 16600
rect 101120 16400 101130 16600
rect 97580 15300 98000 15600
rect 101180 15500 101300 17120
rect 101500 140520 101600 141800
rect 101650 141200 101660 141400
rect 101860 141200 101870 141400
rect 101500 17120 101660 140520
rect 101500 16606 101600 17120
rect 101496 16398 101506 16606
rect 101860 16398 101870 16606
rect 101500 15800 101600 16398
rect 102000 15780 103000 142200
rect 104510 141200 104520 141400
rect 104510 16400 104520 16600
rect 104720 15800 104900 141800
rect 101100 15400 101300 15500
rect 101100 15300 101200 15400
rect 101300 15300 101310 15400
rect 60100 14900 94400 15100
<< via1 >>
rect 58200 143400 59200 144400
rect 68400 143400 69600 144400
rect 75600 143400 76600 144400
rect 82800 143400 84000 144400
rect 90000 143400 91200 144400
rect 97200 143400 98400 144400
rect 63000 142200 64000 143000
rect 40400 133000 42200 133800
rect 41200 129800 41600 130200
rect 48680 131110 48840 131170
rect 49050 131110 49230 131170
rect 49430 131120 49610 131180
rect 49810 131120 49990 131180
rect 50190 131110 50370 131170
rect 50570 131110 50750 131170
rect 48610 130900 48670 131000
rect 48180 130360 48420 130600
rect 48840 130900 48900 131000
rect 48990 130900 49050 131000
rect 49210 130900 49280 131000
rect 49370 130900 49440 131000
rect 49590 130900 49660 131000
rect 49750 130900 49820 131000
rect 49970 130900 50040 131000
rect 50140 130900 50210 131000
rect 50350 130900 50420 131000
rect 50510 130900 50580 131000
rect 48670 130740 48850 130800
rect 48670 128770 48850 128830
rect 48600 128550 48670 128650
rect 49050 130740 49230 130800
rect 49430 130750 49610 130810
rect 49810 130750 49990 130810
rect 50190 130740 50370 130800
rect 48970 130360 49070 130460
rect 49250 130240 49310 130300
rect 49050 130000 49220 130070
rect 49670 130230 49740 130300
rect 50350 130370 50450 130470
rect 50110 130240 50170 130300
rect 50190 130000 50360 130070
rect 49050 128770 49230 128830
rect 49430 128770 49610 128830
rect 49810 128770 49990 128830
rect 50190 128770 50370 128830
rect 50740 130900 50810 131000
rect 50570 130740 50750 130800
rect 50570 128770 50750 128830
rect 48830 128560 48900 128660
rect 49000 128560 49070 128660
rect 49210 128560 49280 128660
rect 49380 128560 49450 128660
rect 49590 128560 49660 128660
rect 49760 128560 49830 128660
rect 49970 128560 50040 128660
rect 50140 128560 50210 128660
rect 50350 128560 50420 128660
rect 50520 128560 50590 128660
rect 51720 130360 51960 130600
rect 51200 130000 51400 130200
rect 50730 128560 50800 128660
rect 48670 128400 48850 128460
rect 49050 128400 49230 128460
rect 49430 128400 49610 128460
rect 49810 128400 49990 128460
rect 50190 128400 50370 128460
rect 50570 128400 50750 128460
rect 48200 116600 48400 116800
rect 43800 112900 44400 113300
rect 43620 111860 43720 112360
rect 43620 92320 43720 92820
rect 44600 111860 44700 112360
rect 45300 112900 45900 113300
rect 45020 111860 45120 112360
rect 44600 92320 44700 92820
rect 45020 92340 45120 92840
rect 46000 111860 46100 112360
rect 48200 113800 48400 114000
rect 46700 112900 47300 113300
rect 48100 112900 48700 113300
rect 46420 111860 46520 112360
rect 46000 92340 46100 92840
rect 46420 92340 46520 92840
rect 47400 111860 47500 112360
rect 47820 111860 47920 112360
rect 47400 92340 47500 92840
rect 47820 92340 47940 92840
rect 48800 111860 48900 112360
rect 49500 112900 50100 113300
rect 49220 111860 49320 112360
rect 48800 92340 48900 92840
rect 47560 91460 47760 91760
rect 49220 92340 49320 92840
rect 50900 112900 51500 113300
rect 50200 111860 50300 112360
rect 50620 111860 50720 112360
rect 50200 92340 50300 92840
rect 50620 92766 50720 92840
rect 50516 92388 50726 92766
rect 50620 92340 50720 92388
rect 51600 111860 51700 112360
rect 51600 92340 51700 92840
rect 46000 90400 46400 90800
rect 43900 87500 44500 87900
rect 43660 86660 43820 87040
rect 43660 66820 43820 67220
rect 44580 86660 44720 87040
rect 44620 66820 44720 67200
rect 47560 88020 47760 88340
rect 45300 87500 45900 87900
rect 45060 86660 45160 87040
rect 45060 66820 45220 67200
rect 46040 86660 46140 87040
rect 45960 66820 46120 67200
rect 46700 87500 47300 87900
rect 48100 87500 48700 87900
rect 46460 86660 46620 87040
rect 46200 66440 46260 66540
rect 46460 66820 46600 67200
rect 47420 86660 47520 87040
rect 47860 86660 48020 87060
rect 47380 66820 47520 67200
rect 47860 66820 48000 67200
rect 48820 86660 48940 87040
rect 49500 87500 50100 87900
rect 48820 66820 48940 67200
rect 49260 86660 49420 87040
rect 49260 66820 49380 67200
rect 49120 66440 49180 66540
rect 50180 86660 50320 87040
rect 50900 87500 51500 87900
rect 50220 66820 50340 67200
rect 50660 86660 50800 87040
rect 50660 66820 50760 67200
rect 51600 86660 51740 87040
rect 51620 66820 51720 67200
rect 45000 51800 45400 52200
rect 46200 54300 46600 54500
rect 47000 54300 47400 54500
rect 46820 51820 46920 52800
rect 47800 54300 48200 54500
rect 47520 49320 47660 50340
rect 48600 54300 49000 54500
rect 48320 50560 48460 51580
rect 49400 54300 49800 54500
rect 49120 49320 49260 50340
rect 50200 54300 50600 54500
rect 49860 51820 49960 52800
rect 45000 37960 45400 38480
rect 51300 37400 51520 37600
rect 50100 37000 50320 37200
rect 49200 35700 49400 35800
rect 52200 35700 52400 35800
rect 49880 35480 49940 35540
rect 50480 35480 50540 35540
rect 51080 35480 51140 35540
rect 51680 35480 51740 35540
rect 49500 35240 49720 35380
rect 50100 35240 50320 35380
rect 50700 35240 50920 35380
rect 51300 35240 51520 35380
rect 51900 35240 52120 35380
rect 49200 34500 49400 34600
rect 52200 34500 52400 34600
rect 49880 34240 49940 34400
rect 50480 34240 50540 34400
rect 51080 34240 51140 34400
rect 51680 34240 51740 34400
rect 49200 33300 49400 33400
rect 52200 33300 52400 33400
rect 49880 33000 49940 33160
rect 50480 33000 50540 33160
rect 51080 33000 51140 33160
rect 51680 33000 51740 33160
rect 49200 32000 49400 32100
rect 52200 32000 52400 32100
rect 49880 31780 49940 31940
rect 50480 31780 50540 31940
rect 51080 31780 51140 31940
rect 51680 31780 51740 31940
rect 49200 30800 49400 30900
rect 52200 30800 52400 30900
rect 49880 30540 49940 30700
rect 50480 30540 50540 30700
rect 51080 30540 51140 30700
rect 51680 30540 51740 30700
rect 49200 29600 49400 29700
rect 52200 29600 52400 29700
rect 49880 29300 49940 29460
rect 50480 29300 50540 29460
rect 51080 29300 51140 29460
rect 51680 29300 51740 29460
rect 49200 28400 49400 28500
rect 52200 28400 52400 28500
rect 49880 28080 49940 28220
rect 50480 28080 50540 28220
rect 51080 28080 51140 28220
rect 51680 28080 51740 28220
rect 49200 27100 49400 27200
rect 52200 27100 52400 27200
rect 49880 26820 49940 26980
rect 50480 26840 50540 27000
rect 51080 26840 51140 27000
rect 51680 26840 51740 27000
rect 49200 25900 49400 26000
rect 52200 25900 52400 26000
rect 49880 25600 49940 25760
rect 50480 25600 50540 25760
rect 51080 25600 51140 25760
rect 51680 25600 51740 25760
rect 49200 24700 49400 24800
rect 52200 24700 52400 24800
rect 49880 24360 49940 24520
rect 50480 24360 50540 24520
rect 51080 24360 51140 24520
rect 51680 24360 51740 24520
rect 49200 23400 49400 23500
rect 52200 23400 52400 23500
rect 49880 23120 49940 23280
rect 50480 23120 50540 23280
rect 51080 23120 51140 23280
rect 51680 23120 51740 23280
rect 49200 22200 49400 22300
rect 49880 21880 49940 22040
rect 50480 21880 50540 22040
rect 51080 21880 51140 22040
rect 52200 22200 52400 22300
rect 51680 21880 51740 22040
rect 49200 20900 49400 21000
rect 52200 20900 52400 21000
rect 49880 20660 49940 20820
rect 50480 20660 50540 20820
rect 51080 20660 51140 20820
rect 51680 20660 51740 20820
rect 49200 19700 49400 19800
rect 52200 19700 52400 19800
rect 49880 19420 49940 19580
rect 50480 19420 50540 19580
rect 51080 19420 51140 19580
rect 51680 19420 51740 19580
rect 49200 18500 49400 18600
rect 52200 18500 52400 18600
rect 49880 18180 49940 18340
rect 50480 18180 50540 18340
rect 51080 18180 51140 18340
rect 51680 18180 51740 18340
rect 49200 17200 49400 17300
rect 52200 17200 52400 17300
rect 49880 17040 49940 17100
rect 50480 17040 50540 17100
rect 51080 17040 51140 17100
rect 51680 17040 51740 17100
rect 49200 15900 49400 16000
rect 52200 15900 52400 16000
rect 51080 15800 51140 15860
rect 62060 141200 62260 141400
rect 62060 16400 62260 16600
rect 66592 142194 67612 142988
rect 70000 142200 71000 143000
rect 74000 142200 75000 143000
rect 77000 142200 78000 143000
rect 81000 142200 82000 143000
rect 85000 142200 86000 143000
rect 88000 142200 89000 143000
rect 92000 142200 93000 143000
rect 95000 142200 96000 143000
rect 99000 142200 100000 143000
rect 102000 142200 103000 143000
rect 64920 141200 65120 141400
rect 64920 16400 65120 16600
rect 65660 141200 65860 141400
rect 65660 16400 65860 16600
rect 68520 141200 68720 141400
rect 68520 16400 68720 16600
rect 69260 141200 69460 141400
rect 69260 16400 69460 16600
rect 72120 141200 72320 141400
rect 72120 16400 72320 16600
rect 72860 141200 73060 141400
rect 72400 15300 72500 15400
rect 72860 16400 73060 16600
rect 75720 141200 75920 141400
rect 75720 16400 75920 16600
rect 76460 141200 76660 141400
rect 76460 16400 76660 16600
rect 79320 141200 79520 141400
rect 79320 16400 79520 16600
rect 80060 141200 80260 141400
rect 79600 15300 79700 15400
rect 80060 16400 80260 16600
rect 82920 141200 83120 141400
rect 82920 16400 83120 16600
rect 83660 141200 83860 141400
rect 83660 16400 83860 16600
rect 86520 141200 86720 141400
rect 86520 16400 86720 16600
rect 87260 141200 87460 141400
rect 86800 15300 86900 15400
rect 87260 16400 87460 16600
rect 90120 141200 90320 141400
rect 90120 16400 90320 16600
rect 90860 141200 91060 141400
rect 90860 16400 91060 16600
rect 93720 141200 93920 141400
rect 93720 16400 93920 16600
rect 94460 141200 94660 141400
rect 94000 15300 94100 15400
rect 94460 16400 94660 16600
rect 97320 141200 97520 141400
rect 97320 16400 97520 16600
rect 98060 141200 98260 141400
rect 98060 16400 98260 16600
rect 100920 141200 101120 141400
rect 100920 16400 101120 16600
rect 101660 141200 101860 141400
rect 101506 16398 101860 16606
rect 104520 141200 104720 141400
rect 104520 16400 104720 16600
rect 101200 15300 101300 15400
<< metal2 >>
rect 38000 144400 98400 145000
rect 38000 143400 58200 144400
rect 59200 143400 68400 144400
rect 69600 143400 75600 144400
rect 76600 143400 82800 144400
rect 84000 143400 90000 144400
rect 91200 143400 97200 144400
rect 38000 140800 40000 143400
rect 58200 143390 59200 143400
rect 68400 143390 69600 143400
rect 75600 143390 76600 143400
rect 82800 143390 84000 143400
rect 90000 143390 91200 143400
rect 97200 143390 98400 143400
rect 63000 143000 64000 143010
rect 70000 143000 71000 143010
rect 74000 143000 75000 143010
rect 77000 143000 78000 143010
rect 81000 143000 82000 143010
rect 85000 143000 86000 143010
rect 88000 143000 89000 143010
rect 92000 143000 93000 143010
rect 95000 143000 96000 143010
rect 99000 143000 100000 143010
rect 102000 143000 103000 143010
rect 38000 139200 38200 140800
rect 39800 139200 40000 140800
rect 38000 139000 40000 139200
rect 59000 142200 63000 143000
rect 64000 142988 70000 143000
rect 64000 142200 66592 142988
rect 40414 134800 52400 134812
rect 52600 134800 54600 134810
rect 40414 133810 52600 134800
rect 40400 133800 52600 133810
rect 42200 133000 52600 133800
rect 40400 132990 52400 133000
rect 40414 132982 52400 132990
rect 49430 131180 49610 131190
rect 47458 131170 47704 131174
rect 48680 131170 48840 131180
rect 49050 131170 49230 131180
rect 47458 131110 48680 131170
rect 48840 131110 49050 131170
rect 49230 131120 49430 131170
rect 49810 131180 49990 131190
rect 49610 131120 49810 131170
rect 50190 131170 50370 131180
rect 50570 131170 50750 131180
rect 49990 131120 50190 131170
rect 49230 131110 50190 131120
rect 50370 131110 50570 131170
rect 47458 131104 48888 131110
rect 41200 130200 41600 130210
rect 47458 130200 47704 131104
rect 48680 131100 48840 131104
rect 49050 131100 49230 131110
rect 50190 131100 50370 131110
rect 50570 131100 50750 131110
rect 48610 131000 48670 131010
rect 48840 131000 48900 131010
rect 48670 130920 48840 130980
rect 48610 130890 48670 130900
rect 48990 131000 49050 131010
rect 48900 130920 48990 130980
rect 48840 130890 48900 130900
rect 49210 131000 49280 131010
rect 49050 130920 49210 130980
rect 48990 130890 49050 130900
rect 49370 131000 49440 131010
rect 49280 130920 49370 130980
rect 49210 130890 49280 130900
rect 49590 131000 49660 131010
rect 49440 130920 49590 130980
rect 49370 130890 49440 130900
rect 49750 131000 49820 131010
rect 49660 130920 49750 130980
rect 49590 130890 49660 130900
rect 49970 131000 50040 131010
rect 49820 130920 49970 130980
rect 49750 130890 49820 130900
rect 50140 131000 50210 131010
rect 50040 130920 50140 130980
rect 49970 130890 50040 130900
rect 50350 131000 50420 131010
rect 50210 130920 50350 130980
rect 50140 130890 50210 130900
rect 50510 131000 50580 131010
rect 50420 130920 50510 130980
rect 50350 130890 50420 130900
rect 50740 131000 50810 131010
rect 50580 130920 50740 130980
rect 50510 130890 50580 130900
rect 50740 130890 50810 130900
rect 49430 130810 49610 130820
rect 48670 130800 48850 130810
rect 49050 130800 49230 130810
rect 48850 130740 49050 130800
rect 49230 130750 49430 130800
rect 49810 130810 49990 130820
rect 49610 130750 49810 130800
rect 50190 130800 50370 130810
rect 50570 130800 50750 130810
rect 49990 130750 50190 130800
rect 49230 130740 50190 130750
rect 50370 130740 50570 130800
rect 48670 130730 48850 130740
rect 49050 130730 49230 130740
rect 50190 130730 50370 130740
rect 50570 130730 50750 130740
rect 48180 130600 48420 130610
rect 51720 130600 51960 130610
rect 48420 130460 49080 130600
rect 48420 130360 48970 130460
rect 49070 130360 49080 130460
rect 50340 130470 51720 130600
rect 50340 130370 50350 130470
rect 50450 130370 51720 130470
rect 50340 130360 51720 130370
rect 48180 130350 48420 130360
rect 48970 130350 49070 130360
rect 51720 130350 51960 130360
rect 49250 130300 49310 130310
rect 49670 130300 49740 130310
rect 50110 130300 50170 130310
rect 49310 130240 49670 130300
rect 49250 130230 49310 130240
rect 49740 130240 50110 130300
rect 50170 130240 52600 130300
rect 50110 130230 50170 130240
rect 49670 130220 49740 130230
rect 41600 130146 47704 130200
rect 51200 130200 51400 130210
rect 41600 130080 47700 130146
rect 41600 130070 49220 130080
rect 41600 130000 49050 130070
rect 41600 129800 47700 130000
rect 49050 129990 49220 130000
rect 50190 130070 51200 130080
rect 50360 130000 51200 130070
rect 52600 130190 54600 130200
rect 50190 129990 50360 130000
rect 51200 129990 51400 130000
rect 41200 129790 41600 129800
rect 48670 128830 48850 128840
rect 49050 128830 49230 128840
rect 49430 128830 49610 128840
rect 49810 128830 49990 128840
rect 50190 128830 50370 128840
rect 50570 128830 50750 128840
rect 48850 128770 49050 128830
rect 49230 128770 49430 128830
rect 49610 128770 49810 128830
rect 49990 128770 50190 128830
rect 50370 128770 50570 128830
rect 48670 128760 48850 128770
rect 49050 128760 49230 128770
rect 49430 128760 49610 128770
rect 49810 128760 49990 128770
rect 50190 128760 50370 128770
rect 50570 128760 50750 128770
rect 48830 128660 48900 128670
rect 49000 128660 49070 128670
rect 49210 128660 49280 128670
rect 49380 128660 49450 128670
rect 49590 128660 49660 128670
rect 49760 128660 49830 128670
rect 49970 128660 50040 128670
rect 50140 128660 50210 128670
rect 50350 128660 50420 128670
rect 50520 128660 50590 128670
rect 50730 128660 50800 128670
rect 48600 128650 48830 128660
rect 48670 128560 48830 128650
rect 48900 128560 49000 128660
rect 49070 128560 49210 128660
rect 49280 128560 49380 128660
rect 49450 128560 49590 128660
rect 49660 128560 49760 128660
rect 49830 128560 49970 128660
rect 50040 128560 50140 128660
rect 50210 128560 50350 128660
rect 50420 128560 50520 128660
rect 50590 128560 50730 128660
rect 48830 128550 48900 128560
rect 49000 128550 49070 128560
rect 49210 128550 49280 128560
rect 49380 128550 49450 128560
rect 49590 128550 49660 128560
rect 49760 128550 49830 128560
rect 49970 128550 50040 128560
rect 50140 128550 50210 128560
rect 50350 128550 50420 128560
rect 50520 128550 50590 128560
rect 50730 128550 50800 128560
rect 48600 128540 48670 128550
rect 48670 128460 50750 128470
rect 48850 128410 49050 128460
rect 48670 128390 48850 128400
rect 49230 128410 49430 128460
rect 49050 128390 49230 128400
rect 49610 128410 49810 128460
rect 49430 128390 49610 128400
rect 49990 128410 50190 128460
rect 49810 128390 49990 128400
rect 50370 128410 50570 128460
rect 50190 128390 50370 128400
rect 50570 128390 50750 128400
rect 48200 116800 48400 116810
rect 48200 114000 48400 116600
rect 48200 113790 48400 113800
rect 36000 113300 36800 113310
rect 43800 113300 44400 113310
rect 45300 113300 45900 113310
rect 46700 113300 47300 113310
rect 48100 113300 48700 113310
rect 49500 113300 50100 113310
rect 50900 113300 51500 113310
rect 36800 112900 43800 113300
rect 44400 112900 45300 113300
rect 45900 112900 46700 113300
rect 47300 112900 48100 113300
rect 48700 112900 49500 113300
rect 50100 113298 50460 113300
rect 50782 113298 50900 113300
rect 50100 112900 50900 113298
rect 51500 112900 51600 113300
rect 36000 112890 36800 112900
rect 43800 112890 44400 112900
rect 45300 112890 45900 112900
rect 46700 112890 47300 112900
rect 48100 112890 48700 112900
rect 49500 112890 50100 112900
rect 50246 112894 51600 112900
rect 50900 112890 51500 112894
rect 43620 112360 43720 112370
rect 44600 112360 44700 112370
rect 43720 111900 44600 112280
rect 43620 111850 43720 111860
rect 45020 112360 45120 112370
rect 44700 112276 44870 112280
rect 44988 112276 45020 112280
rect 44700 111902 45020 112276
rect 44700 111900 44870 111902
rect 44988 111900 45020 111902
rect 44600 111850 44700 111860
rect 46000 112360 46100 112370
rect 45120 111900 46000 112280
rect 45020 111850 45120 111860
rect 46420 112360 46520 112370
rect 46100 111900 46420 112280
rect 46000 111850 46100 111860
rect 47400 112360 47500 112370
rect 46520 111900 47400 112280
rect 46420 111850 46520 111860
rect 47820 112360 47920 112370
rect 47500 111900 47820 112280
rect 47400 111850 47500 111860
rect 48800 112360 48900 112370
rect 47920 111900 48800 112280
rect 47820 111850 47920 111860
rect 49220 112360 49320 112370
rect 48900 111900 49220 112280
rect 48800 111850 48900 111860
rect 50200 112360 50300 112370
rect 49320 111900 50200 112280
rect 49220 111850 49320 111860
rect 50620 112360 50720 112370
rect 50300 111900 50620 112280
rect 50200 111850 50300 111860
rect 51600 112360 51700 112370
rect 50720 111900 51600 112280
rect 50620 111850 50720 111860
rect 51600 111850 51700 111860
rect 59000 105400 59400 142200
rect 63000 142190 64000 142200
rect 67612 142200 70000 142988
rect 71000 142200 74000 143000
rect 75000 142200 77000 143000
rect 78000 142200 81000 143000
rect 82000 142200 85000 143000
rect 86000 142200 88000 143000
rect 89000 142200 92000 143000
rect 93000 142200 95000 143000
rect 96000 142200 99000 143000
rect 100000 142200 102000 143000
rect 66592 142184 67612 142194
rect 70000 142190 71000 142200
rect 74000 142190 75000 142200
rect 77000 142190 78000 142200
rect 81000 142190 82000 142200
rect 85000 142190 86000 142200
rect 88000 142190 89000 142200
rect 92000 142190 93000 142200
rect 95000 142190 96000 142200
rect 99000 142190 100000 142200
rect 102000 142190 103000 142200
rect 62060 141400 62260 141410
rect 64920 141400 65120 141410
rect 65660 141400 65860 141410
rect 68520 141400 68720 141410
rect 69260 141400 69460 141410
rect 72120 141400 72320 141410
rect 72860 141400 73060 141410
rect 75720 141400 75920 141410
rect 76460 141400 76660 141410
rect 79320 141400 79520 141410
rect 80060 141400 80260 141410
rect 82920 141400 83120 141410
rect 83660 141400 83860 141410
rect 86520 141400 86720 141410
rect 87260 141400 87460 141410
rect 90120 141400 90320 141410
rect 90860 141400 91060 141410
rect 93720 141400 93920 141410
rect 94460 141400 94660 141410
rect 97320 141400 97520 141410
rect 98060 141400 98260 141410
rect 100920 141400 101120 141410
rect 101660 141400 101860 141410
rect 104520 141400 104720 141410
rect 62000 141200 62060 141400
rect 62260 141200 64920 141400
rect 65120 141200 65660 141400
rect 65860 141200 68520 141400
rect 68720 141200 69260 141400
rect 69460 141200 72120 141400
rect 72320 141200 72860 141400
rect 73060 141200 75720 141400
rect 75920 141200 76460 141400
rect 76660 141200 79320 141400
rect 79520 141200 80060 141400
rect 80260 141200 82920 141400
rect 83120 141200 83660 141400
rect 83860 141200 86520 141400
rect 86720 141200 87260 141400
rect 87460 141200 90120 141400
rect 90320 141200 90860 141400
rect 91060 141200 93720 141400
rect 93920 141200 94460 141400
rect 94660 141200 97320 141400
rect 97520 141200 98060 141400
rect 98260 141200 100920 141400
rect 101120 141200 101660 141400
rect 101860 141200 104520 141400
rect 104720 141200 104800 141400
rect 62060 141190 62260 141200
rect 64920 141190 65120 141200
rect 65660 141190 65860 141200
rect 68520 141190 68720 141200
rect 69260 141190 69460 141200
rect 72120 141190 72320 141200
rect 72860 141190 73060 141200
rect 75720 141190 75920 141200
rect 76460 141190 76660 141200
rect 79320 141190 79520 141200
rect 80060 141190 80260 141200
rect 82920 141190 83120 141200
rect 83660 141190 83860 141200
rect 86520 141190 86720 141200
rect 87260 141190 87460 141200
rect 90120 141190 90320 141200
rect 90860 141190 91060 141200
rect 93720 141190 93920 141200
rect 94460 141190 94660 141200
rect 97320 141190 97520 141200
rect 98060 141190 98260 141200
rect 100920 141190 101120 141200
rect 101660 141190 101860 141200
rect 104520 141190 104720 141200
rect 53200 105000 59400 105400
rect 45020 92840 45120 92850
rect 43620 92820 43720 92830
rect 44600 92820 44700 92830
rect 43720 92380 44600 92760
rect 43620 92310 43720 92320
rect 44700 92382 45020 92760
rect 44700 92380 44854 92382
rect 44986 92380 45020 92382
rect 46000 92840 46100 92850
rect 45120 92380 46000 92760
rect 45020 92330 45120 92340
rect 46420 92840 46520 92850
rect 46100 92380 46420 92760
rect 46000 92330 46100 92340
rect 47400 92840 47500 92850
rect 46520 92380 47400 92760
rect 46420 92330 46520 92340
rect 47820 92840 47940 92850
rect 47500 92380 47820 92760
rect 47400 92330 47500 92340
rect 48800 92840 48900 92850
rect 47940 92380 48800 92760
rect 47820 92330 47940 92340
rect 49220 92840 49320 92850
rect 48900 92380 49220 92760
rect 48800 92330 48900 92340
rect 50200 92840 50300 92850
rect 49320 92380 50200 92760
rect 49220 92330 49320 92340
rect 50620 92840 50720 92850
rect 50516 92766 50620 92776
rect 51600 92840 51700 92850
rect 50720 92766 50726 92776
rect 50300 92388 50516 92760
rect 50726 92388 51600 92760
rect 50300 92380 50620 92388
rect 50516 92378 50620 92380
rect 50200 92330 50300 92340
rect 50720 92380 51600 92388
rect 50720 92378 50726 92380
rect 50620 92330 50720 92340
rect 51600 92330 51700 92340
rect 44600 92310 44700 92320
rect 47560 91760 47760 91770
rect 47560 90956 47760 91460
rect 47558 90908 47760 90956
rect 36000 90800 36800 90810
rect 46000 90800 46400 90810
rect 36800 90400 46000 90800
rect 47558 90562 47756 90908
rect 47558 90510 47760 90562
rect 36000 90390 36800 90400
rect 46000 90390 46400 90400
rect 47560 90200 47760 90510
rect 53200 90200 53600 105000
rect 47560 89800 53600 90200
rect 47560 88340 47760 89800
rect 47560 88010 47760 88020
rect 36000 87900 36800 87910
rect 43900 87900 44500 87910
rect 45300 87900 45900 87910
rect 46700 87900 47300 87910
rect 48100 87900 48700 87910
rect 49500 87900 50100 87910
rect 50900 87900 51500 87910
rect 36800 87500 43900 87900
rect 44500 87500 45300 87900
rect 45900 87500 46700 87900
rect 47300 87500 48100 87900
rect 48700 87500 49500 87900
rect 50100 87500 50900 87900
rect 51500 87500 52000 87900
rect 36000 87490 36800 87500
rect 43900 87490 44500 87500
rect 45300 87490 45900 87500
rect 46700 87490 47300 87500
rect 48100 87490 48700 87500
rect 49500 87490 50100 87500
rect 50900 87490 51500 87500
rect 47860 87060 48020 87070
rect 43660 87040 43820 87050
rect 44580 87040 44720 87050
rect 45060 87040 45160 87050
rect 46040 87040 46140 87050
rect 46460 87040 46620 87050
rect 47420 87040 47520 87050
rect 43820 86660 44580 87040
rect 44720 86660 45060 87040
rect 45160 86660 46040 87040
rect 46140 86660 46460 87040
rect 46620 86660 47420 87040
rect 47520 86660 47860 87040
rect 48820 87040 48940 87050
rect 49260 87040 49420 87050
rect 50180 87040 50320 87050
rect 50660 87040 50800 87050
rect 51600 87040 51740 87050
rect 48020 86660 48820 87040
rect 48940 86660 49260 87040
rect 49420 86660 50180 87040
rect 50320 86660 50660 87040
rect 50800 86660 51600 87040
rect 43660 86650 43820 86660
rect 44580 86650 44720 86660
rect 45060 86650 45160 86660
rect 46040 86650 46140 86660
rect 46460 86650 46620 86660
rect 47420 86650 47520 86660
rect 47860 86650 48020 86660
rect 48820 86650 48940 86660
rect 49260 86650 49420 86660
rect 50180 86650 50320 86660
rect 50660 86650 50800 86660
rect 51600 86650 51740 86660
rect 43660 67220 43820 67230
rect 44620 67200 44720 67210
rect 45060 67200 45220 67210
rect 45960 67200 46120 67210
rect 46460 67200 46600 67210
rect 47380 67200 47520 67210
rect 47860 67200 48000 67210
rect 48820 67200 48940 67210
rect 49260 67200 49380 67210
rect 50220 67200 50340 67210
rect 50660 67200 50760 67210
rect 51620 67200 51720 67210
rect 43820 66820 44620 67200
rect 44720 66820 45060 67200
rect 45220 66820 45960 67200
rect 46120 66820 46460 67200
rect 46600 66820 47380 67200
rect 47520 66820 47860 67200
rect 48000 66820 48820 67200
rect 48940 66820 49260 67200
rect 49380 66820 50220 67200
rect 50340 66820 50660 67200
rect 50760 66820 51620 67200
rect 43660 66810 43820 66820
rect 44620 66810 44720 66820
rect 45060 66810 45220 66820
rect 45960 66810 46120 66820
rect 46460 66810 46600 66820
rect 47380 66810 47520 66820
rect 47860 66810 48000 66820
rect 48820 66810 48940 66820
rect 49260 66810 49380 66820
rect 50220 66810 50340 66820
rect 50660 66810 50760 66820
rect 51620 66810 51720 66820
rect 46200 66540 46260 66550
rect 46200 65400 46260 66440
rect 49120 66540 49180 66550
rect 49120 65400 49180 66440
rect 46200 65000 59800 65400
rect 36000 54600 36800 54610
rect 36800 54500 54200 54600
rect 36800 54300 46200 54500
rect 46600 54300 47000 54500
rect 47400 54300 47800 54500
rect 48200 54300 48600 54500
rect 49000 54300 49400 54500
rect 49800 54300 50200 54500
rect 50600 54300 54200 54500
rect 36000 54290 36800 54300
rect 46200 54290 46600 54300
rect 47000 54290 47400 54300
rect 47800 54290 48200 54300
rect 48600 54290 49000 54300
rect 49400 54290 49800 54300
rect 50200 54290 50600 54300
rect 46820 52800 46920 52810
rect 45000 52200 45400 52210
rect 45400 51820 46820 52200
rect 49860 52800 49960 52810
rect 46920 51820 49860 52200
rect 49960 51820 50000 52200
rect 45400 51800 50000 51820
rect 45000 51790 45400 51800
rect 48320 51580 48460 51590
rect 46020 50560 48320 50900
rect 54000 50900 54200 54300
rect 48460 50560 54220 50900
rect 48320 50550 48460 50560
rect 47520 50340 47660 50350
rect 38000 49800 40000 49810
rect 40000 49660 40600 49800
rect 40000 49320 47520 49660
rect 49120 50340 49260 50350
rect 47660 49320 49120 49660
rect 40000 49200 40600 49320
rect 47520 49310 47660 49320
rect 49120 49310 49260 49320
rect 38000 49190 40000 49200
rect 45000 38480 45400 38490
rect 45400 37960 52120 38480
rect 45000 37950 45400 37960
rect 49200 35800 49400 35810
rect 49200 34600 49400 35700
rect 49500 35380 49720 37960
rect 50100 37200 50320 37210
rect 49500 35230 49720 35240
rect 49880 35540 49940 35550
rect 49200 33400 49400 34500
rect 49200 32100 49400 33300
rect 49200 30900 49400 32000
rect 49200 29700 49400 30800
rect 49200 28500 49400 29600
rect 49200 27200 49400 28400
rect 49200 26000 49400 27100
rect 49200 24800 49400 25900
rect 49200 23500 49400 24700
rect 49200 22300 49400 23400
rect 49200 21000 49400 22200
rect 49200 19800 49400 20900
rect 36000 19200 36800 19210
rect 36800 18800 44200 19200
rect 36000 18790 36800 18800
rect 43800 15600 44200 18800
rect 49200 18600 49400 19700
rect 49200 17300 49400 18500
rect 49200 16000 49400 17200
rect 49200 15890 49400 15900
rect 49880 34400 49940 35480
rect 50100 35380 50320 37000
rect 50100 35230 50320 35240
rect 50480 35540 50540 35550
rect 49880 33160 49940 34240
rect 49880 31940 49940 33000
rect 49880 30700 49940 31780
rect 49880 29460 49940 30540
rect 49880 28220 49940 29300
rect 49880 26980 49940 28080
rect 49880 25760 49940 26820
rect 49880 24520 49940 25600
rect 49880 23280 49940 24360
rect 49880 22040 49940 23120
rect 49880 20820 49940 21880
rect 49880 19580 49940 20660
rect 49880 18340 49940 19420
rect 49880 17100 49940 18180
rect 49880 15700 49940 17040
rect 50480 34400 50540 35480
rect 50700 35380 50920 37960
rect 51300 37600 51520 37610
rect 50700 35230 50920 35240
rect 51080 35540 51140 35550
rect 50480 33160 50540 34240
rect 50480 31940 50540 33000
rect 50480 30700 50540 31780
rect 50480 29460 50540 30540
rect 50480 28220 50540 29300
rect 50480 27000 50540 28080
rect 50480 25760 50540 26840
rect 50480 24520 50540 25600
rect 50480 23280 50540 24360
rect 50480 22040 50540 23120
rect 50480 20820 50540 21880
rect 50480 19580 50540 20660
rect 50480 18340 50540 19420
rect 50480 17100 50540 18180
rect 50480 15700 50540 17040
rect 49880 15600 50540 15700
rect 43800 15200 50540 15600
rect 51080 34400 51140 35480
rect 51300 35380 51520 37400
rect 51300 35230 51520 35240
rect 51680 35540 51740 35550
rect 51080 33160 51140 34240
rect 51080 31940 51140 33000
rect 51080 30700 51140 31780
rect 51080 29460 51140 30540
rect 51080 28220 51140 29300
rect 51080 27000 51140 28080
rect 51080 25760 51140 26840
rect 51080 24520 51140 25600
rect 51080 23280 51140 24360
rect 51080 22040 51140 23120
rect 51080 20820 51140 21880
rect 51080 19580 51140 20660
rect 51080 18340 51140 19420
rect 51080 17100 51140 18180
rect 51080 15860 51140 17040
rect 51080 15700 51140 15800
rect 51680 34400 51740 35480
rect 51900 35380 52120 37960
rect 51900 35230 52120 35240
rect 52200 35800 52400 35810
rect 51680 33160 51740 34240
rect 51680 31940 51740 33000
rect 51680 30700 51740 31780
rect 51680 29460 51740 30540
rect 51680 28220 51740 29300
rect 51680 27000 51740 28080
rect 51680 25760 51740 26840
rect 51680 24520 51740 25600
rect 51680 23280 51740 24360
rect 51680 22040 51740 23120
rect 51680 20820 51740 21880
rect 51680 19580 51740 20660
rect 51680 18340 51740 19420
rect 51680 17100 51740 18180
rect 51680 15700 51740 17040
rect 52200 34600 52400 35700
rect 52200 33400 52400 34500
rect 52200 32100 52400 33300
rect 52200 30900 52400 32000
rect 52200 29700 52400 30800
rect 52200 28500 52400 29600
rect 52200 27200 52400 28400
rect 52200 26000 52400 27100
rect 52200 24800 52400 25900
rect 52200 23500 52400 24700
rect 52200 22300 52400 23400
rect 52200 21000 52400 22200
rect 52200 19800 52400 20900
rect 52200 18600 52400 19700
rect 52200 17300 52400 18500
rect 52200 16000 52400 17200
rect 52200 15890 52400 15900
rect 36000 14800 36800 14810
rect 51080 14800 51740 15700
rect 59400 15400 59800 65000
rect 62060 16600 62260 16610
rect 64920 16600 65120 16610
rect 65660 16600 65860 16610
rect 68520 16600 68720 16610
rect 69260 16600 69460 16610
rect 72120 16600 72320 16610
rect 72860 16600 73060 16610
rect 75720 16600 75920 16610
rect 76460 16600 76660 16610
rect 79320 16600 79520 16610
rect 80060 16600 80260 16610
rect 82920 16600 83120 16610
rect 83660 16600 83860 16610
rect 86520 16600 86720 16610
rect 87260 16600 87460 16610
rect 90120 16600 90320 16610
rect 90860 16600 91060 16610
rect 93720 16600 93920 16610
rect 94460 16600 94660 16610
rect 97320 16600 97520 16610
rect 98060 16600 98260 16610
rect 100920 16600 101120 16610
rect 101506 16606 101860 16616
rect 62000 16400 62060 16600
rect 62260 16400 64920 16600
rect 65120 16400 65660 16600
rect 65860 16400 68520 16600
rect 68720 16400 69260 16600
rect 69460 16400 72120 16600
rect 72320 16400 72860 16600
rect 73060 16400 75720 16600
rect 75920 16400 76460 16600
rect 76660 16400 79320 16600
rect 79520 16400 80060 16600
rect 80260 16400 82920 16600
rect 83120 16400 83660 16600
rect 83860 16400 86520 16600
rect 86720 16400 87260 16600
rect 87460 16400 90120 16600
rect 90320 16400 90860 16600
rect 91060 16400 93720 16600
rect 93920 16400 94460 16600
rect 94660 16400 97320 16600
rect 97520 16400 98060 16600
rect 98260 16400 100920 16600
rect 101120 16400 101506 16600
rect 62060 16390 62260 16400
rect 64920 16390 65120 16400
rect 65660 16390 65860 16400
rect 68520 16390 68720 16400
rect 69260 16390 69460 16400
rect 72120 16390 72320 16400
rect 72860 16390 73060 16400
rect 75720 16390 75920 16400
rect 76460 16390 76660 16400
rect 79320 16390 79520 16400
rect 80060 16390 80260 16400
rect 82920 16390 83120 16400
rect 83660 16390 83860 16400
rect 86520 16390 86720 16400
rect 87260 16390 87460 16400
rect 90120 16390 90320 16400
rect 90860 16390 91060 16400
rect 93720 16390 93920 16400
rect 94460 16390 94660 16400
rect 97320 16390 97520 16400
rect 98060 16390 98260 16400
rect 100920 16390 101120 16400
rect 104520 16600 104720 16610
rect 101860 16400 104520 16600
rect 104720 16400 104800 16600
rect 101506 16388 101860 16398
rect 104520 16390 104720 16400
rect 72400 15400 72500 15410
rect 79600 15400 79700 15410
rect 86800 15400 86900 15410
rect 94000 15400 94100 15410
rect 101200 15400 101300 15410
rect 59400 15300 72400 15400
rect 72500 15300 79600 15400
rect 79700 15300 86800 15400
rect 86900 15300 94000 15400
rect 94100 15300 101200 15400
rect 101300 15300 101400 15400
rect 59400 15200 101400 15300
rect 36800 14400 51740 14800
rect 36000 14390 36800 14400
<< via2 >>
rect 38200 139200 39800 140800
rect 52600 130200 54600 134800
rect 36000 112900 36800 113300
rect 36000 90400 36800 90800
rect 36000 87500 36800 87900
rect 36000 54300 36800 54600
rect 38000 49200 40000 49800
rect 36000 18800 36800 19200
rect 36000 14400 36800 14800
<< metal3 >>
rect 32800 143000 54600 145000
rect 32800 140800 40000 141000
rect 32800 139200 38200 140800
rect 39800 139200 40000 140800
rect 32800 139000 40000 139200
rect 32800 113400 36000 114000
rect 32800 113305 36800 113400
rect 32800 113300 36810 113305
rect 32800 112900 36000 113300
rect 36800 112900 36810 113300
rect 32800 112895 36810 112900
rect 32800 112800 36800 112895
rect 32800 112000 36000 112800
rect 32800 91000 36000 92000
rect 32800 90805 36800 91000
rect 32800 90800 36810 90805
rect 32800 90400 36000 90800
rect 36800 90400 36810 90800
rect 32800 90395 36810 90400
rect 32800 90200 36800 90395
rect 32800 90000 36000 90200
rect 32800 87905 36800 88000
rect 32800 87900 36810 87905
rect 32800 87500 36000 87900
rect 36800 87500 36810 87900
rect 32800 87495 36810 87500
rect 32800 87400 36800 87495
rect 32800 86000 36000 87400
rect 32800 54700 36000 56000
rect 32800 54605 36800 54700
rect 32800 54600 36810 54605
rect 32800 54300 36000 54600
rect 36800 54300 36810 54600
rect 32800 54295 36810 54300
rect 32800 54200 36800 54295
rect 32800 54000 36000 54200
rect 38000 49805 40000 139000
rect 52600 134805 54600 143000
rect 52590 134800 54610 134805
rect 52590 130200 52600 134800
rect 54600 130200 54610 134800
rect 52590 130195 54610 130200
rect 37990 49800 40010 49805
rect 37990 49200 38000 49800
rect 40000 49200 40010 49800
rect 37990 49195 40010 49200
rect 32800 19205 36000 20000
rect 32800 19200 36810 19205
rect 32800 18800 36000 19200
rect 36800 18800 36810 19200
rect 32800 18795 36810 18800
rect 32800 18000 36000 18795
rect 32800 14805 36000 16000
rect 32800 14800 36810 14805
rect 32800 14400 36000 14800
rect 36800 14400 36810 14800
rect 32800 14395 36810 14400
rect 32800 14000 36000 14395
use sky130_fd_pr__nfet_01v8_3ZAA45  sky130_fd_pr__nfet_01v8_3ZAA45_0
timestamp 1695666882
transform 1 0 50278 0 1 129458
box -158 -588 158 588
use sky130_fd_pr__nfet_01v8_AH5E2K  sky130_fd_pr__nfet_01v8_AH5E2K_0
timestamp 1695666081
transform 1 0 49758 0 1 112078
box -558 -588 558 588
use sky130_fd_pr__nfet_01v8_MHE452  sky130_fd_pr__nfet_01v8_MHE452_0
timestamp 1695666882
transform 1 0 48758 0 1 129783
box -158 -1383 158 1383
use sky130_fd_pr__nfet_01v8_QP5WRD  sky130_fd_pr__nfet_01v8_QP5WRD_0
timestamp 1695666081
transform 1 0 46958 0 1 102334
box -558 -9114 558 9114
use sky130_fd_pr__nfet_01v8_SCE452  sky130_fd_pr__nfet_01v8_SCE452_0
timestamp 1695666882
transform 1 0 49518 0 1 130963
box -158 -213 158 213
use sky130_fd_pr__nfet_01v8_SCE452  sky130_fd_pr__nfet_01v8_SCE452_1
timestamp 1695666882
transform 1 0 49518 0 1 128613
box -158 -213 158 213
use sky130_fd_pr__nfet_01v8_SCE452  sky130_fd_pr__nfet_01v8_SCE452_2
timestamp 1695666882
transform 1 0 49138 0 1 128613
box -158 -213 158 213
use sky130_fd_pr__nfet_01v8_SCE452  sky130_fd_pr__nfet_01v8_SCE452_3
timestamp 1695666882
transform 1 0 49898 0 1 129553
box -158 -213 158 213
use sky130_fd_pr__nfet_01v8_VT3ZQW  sky130_fd_pr__nfet_01v8_VT3ZQW_0
timestamp 1695667127
transform 1 0 50278 0 1 130953
box -158 -213 158 213
use sky130_fd_pr__nfet_01v8_WK8VRD  sky130_fd_pr__nfet_01v8_WK8VRD_0
timestamp 1695666081
transform 1 0 51158 0 1 102332
box -558 -10332 558 10332
use sky130_fd_pr__pfet_01v8_7DHACV  sky130_fd_pr__pfet_01v8_7DHACV_0
timestamp 1695664993
transform 1 0 51112 0 1 26292
box -112 -9252 112 9252
use sky130_fd_pr__pfet_01v8_8DHNHY  sky130_fd_pr__pfet_01v8_8DHNHY_0
timestamp 1695664993
transform 1 0 52312 0 1 26288
box -112 -10488 112 10488
use sky130_fd_pr__pfet_01v8_C2U9V5  sky130_fd_pr__pfet_01v8_C2U9V5_0
timestamp 1695665377
transform 1 0 49594 0 1 48600
box -394 -600 394 600
use sky130_fd_pr__pfet_01v8_E769TZ  sky130_fd_pr__pfet_01v8_E769TZ_0
timestamp 1695663670
transform 1 0 103194 0 1 78818
box -1594 -63018 1594 63018
use sky130_fd_pr__pfet_01v8_F76D73  sky130_fd_pr__pfet_01v8_F76D73_0
timestamp 1695663670
transform 1 0 95994 0 1 78822
box -1594 -61782 1594 61782
use sky130_fd_pr__pfet_01v8_MGA63L  sky130_fd_pr__pfet_01v8_MGA63L_0
timestamp 1695664993
transform 1 0 51712 0 1 36180
box -112 -600 112 600
use sky130_fd_pr__pfet_01v8_P2UXFR  sky130_fd_pr__pfet_01v8_P2UXFR_0
timestamp 1695665377
transform 1 0 47994 0 1 50458
box -394 -1218 394 1218
use sky130_fd_pr__pfet_01v8_RRU5GE  sky130_fd_pr__pfet_01v8_RRU5GE_0
timestamp 1695665377
transform 1 0 47194 0 1 51076
box -394 -1836 394 1836
use sky130_fd_pr__pfet_01v8_RRUZAE  sky130_fd_pr__pfet_01v8_RRUZAE_0
timestamp 1695665377
transform 1 0 50394 0 1 51072
box -394 -3072 394 3072
use sky130_fd_pr__pfet_01v8_SKU9VM  sky130_fd_pr__pfet_01v8_SKU9VM_0
timestamp 1695665689
transform 1 0 45594 0 1 86780
box -594 -600 594 600
use sky130_fd_pr__pfet_01v8_UDM5A5  sky130_fd_pr__pfet_01v8_UDM5A5_0
timestamp 1695665689
transform 1 0 49794 0 1 76892
box -594 -9252 594 9252
use sky130_fd_pr__pfet_01v8_UDMRD5  sky130_fd_pr__pfet_01v8_UDMRD5_0
timestamp 1695665689
transform 1 0 51194 0 1 76888
box -594 -10488 594 10488
use sky130_fd_pr__pfet_01v8_ZLZ7XS  sky130_fd_pr__pfet_01v8_ZLZ7XS_0
timestamp 1695663670
transform 1 0 99594 0 1 141240
box -1594 -600 1594 600
use sky130_fd_pr__pfet_01v8_F76D73  XM1_1
timestamp 1695663670
transform 1 0 74394 0 1 78822
box -1594 -61782 1594 61782
use sky130_fd_pr__pfet_01v8_F76D73  XM1_2
timestamp 1695663670
transform 1 0 81594 0 1 78822
box -1594 -61782 1594 61782
use sky130_fd_pr__pfet_01v8_F76D73  XM1_3
timestamp 1695663670
transform 1 0 88794 0 1 78822
box -1594 -61782 1594 61782
use sky130_fd_pr__pfet_01v8_F76D73  XM1
timestamp 1695663670
transform 1 0 67194 0 1 78822
box -1594 -61782 1594 61782
use sky130_fd_pr__pfet_01v8_UDM5A5  XM2_1
timestamp 1695665689
transform 1 0 48394 0 1 76892
box -594 -9252 594 9252
use sky130_fd_pr__pfet_01v8_UDMRD5  XM2_dummy_2
timestamp 1695665689
transform 1 0 44194 0 1 76888
box -594 -10488 594 10488
use sky130_fd_pr__pfet_01v8_SKU9VM  XM2_dummy_3
timestamp 1695665689
transform 1 0 45594 0 1 67000
box -594 -600 594 600
use sky130_fd_pr__pfet_01v8_SKU9VM  XM2_dummy_4
timestamp 1695665689
transform 1 0 46994 0 1 67000
box -594 -600 594 600
use sky130_fd_pr__pfet_01v8_SKU9VM  XM2_dummy_5
timestamp 1695665689
transform 1 0 48394 0 1 67000
box -594 -600 594 600
use sky130_fd_pr__pfet_01v8_SKU9VM  XM2_dummy_6
timestamp 1695665689
transform 1 0 49794 0 1 67000
box -594 -600 594 600
use sky130_fd_pr__pfet_01v8_SKU9VM  XM2_dummy_7
timestamp 1695665689
transform 1 0 46994 0 1 86780
box -594 -600 594 600
use sky130_fd_pr__pfet_01v8_SKU9VM  XM2_dummy_9
timestamp 1695665689
transform 1 0 49794 0 1 86780
box -594 -600 594 600
use sky130_fd_pr__pfet_01v8_SKU9VM  XM2_dummy_10
timestamp 1695665689
transform 1 0 48394 0 1 86780
box -594 -600 594 600
use sky130_fd_pr__pfet_01v8_UDM5A5  XM2
timestamp 1695665689
transform 1 0 46994 0 1 76892
box -594 -9252 594 9252
use sky130_fd_pr__nfet_01v8_WK8VRD  XM3_dummy_1
timestamp 1695666081
transform 1 0 44158 0 1 102332
box -558 -10332 558 10332
use sky130_fd_pr__nfet_01v8_AH5E2K  XM3_dummy_3
timestamp 1695666081
transform 1 0 46958 0 1 112078
box -558 -588 558 588
use sky130_fd_pr__nfet_01v8_AH5E2K  XM3_dummy_4
timestamp 1695666081
transform 1 0 48358 0 1 112078
box -558 -588 558 588
use sky130_fd_pr__nfet_01v8_AH5E2K  XM3_dummy_6
timestamp 1695666081
transform 1 0 45558 0 1 112078
box -558 -588 558 588
use sky130_fd_pr__nfet_01v8_AH5E2K  XM3_dummy_7
timestamp 1695666081
transform 1 0 49758 0 1 92588
box -558 -588 558 588
use sky130_fd_pr__nfet_01v8_AH5E2K  XM3_dummy_8
timestamp 1695666081
transform 1 0 46958 0 1 92588
box -558 -588 558 588
use sky130_fd_pr__nfet_01v8_AH5E2K  XM3_dummy_9
timestamp 1695666081
transform 1 0 45558 0 1 92588
box -558 -588 558 588
use sky130_fd_pr__nfet_01v8_AH5E2K  XM3_dummy_10
timestamp 1695666081
transform 1 0 48358 0 1 92588
box -558 -588 558 588
use sky130_fd_pr__nfet_01v8_QP5WRD  XM3
timestamp 1695666081
transform 1 0 48358 0 1 102334
box -558 -9114 558 9114
use sky130_fd_pr__nfet_01v8_MHE452  XM4_dummy_2
timestamp 1695666882
transform 1 0 50658 0 1 129783
box -158 -1383 158 1383
use sky130_fd_pr__nfet_01v8_SCE452  XM4_dummy_3
timestamp 1695666882
transform 1 0 50278 0 1 128613
box -158 -213 158 213
use sky130_fd_pr__nfet_01v8_SCE452  XM4_dummy_7
timestamp 1695666882
transform 1 0 49898 0 1 128613
box -158 -213 158 213
use sky130_fd_pr__nfet_01v8_SCE452  XM4_dummy_9
timestamp 1695666882
transform 1 0 49138 0 1 130953
box -158 -213 158 213
use sky130_fd_pr__nfet_01v8_SCE452  XM4_dummy_10
timestamp 1695666882
transform 1 0 49898 0 1 130963
box -158 -213 158 213
use sky130_fd_pr__nfet_01v8_3ZAA45  XM4
timestamp 1695666882
transform 1 0 49138 0 1 129458
box -158 -588 158 588
use sky130_fd_pr__pfet_01v8_7DHACV  XM5_1
timestamp 1695664993
transform 1 0 50512 0 1 26292
box -112 -9252 112 9252
use sky130_fd_pr__pfet_01v8_8DHNHY  XM5_dummy_1
timestamp 1695664993
transform 1 0 49312 0 1 26288
box -112 -10488 112 10488
use sky130_fd_pr__pfet_01v8_MGA63L  XM5_dummy_3
timestamp 1695664993
transform 1 0 49912 0 1 16400
box -112 -600 112 600
use sky130_fd_pr__pfet_01v8_MGA63L  XM5_dummy_4
timestamp 1695664993
transform 1 0 50512 0 1 16400
box -112 -600 112 600
use sky130_fd_pr__pfet_01v8_MGA63L  XM5_dummy_5
timestamp 1695664993
transform 1 0 51112 0 1 16400
box -112 -600 112 600
use sky130_fd_pr__pfet_01v8_MGA63L  XM5_dummy_6
timestamp 1695664993
transform 1 0 51112 0 1 36180
box -112 -600 112 600
use sky130_fd_pr__pfet_01v8_MGA63L  XM5_dummy_7
timestamp 1695664993
transform 1 0 51712 0 1 16400
box -112 -600 112 600
use sky130_fd_pr__pfet_01v8_MGA63L  XM5_dummy_8
timestamp 1695664993
transform 1 0 49912 0 1 36180
box -112 -600 112 600
use sky130_fd_pr__pfet_01v8_MGA63L  XM5_dummy_10
timestamp 1695664993
transform 1 0 50512 0 1 36180
box -112 -600 112 600
use sky130_fd_pr__pfet_01v8_7DHACV  XM5
timestamp 1695664993
transform 1 0 49912 0 1 26292
box -112 -9252 112 9252
use sky130_fd_pr__nfet_01v8_VT3ZQW  XM6_1
timestamp 1695667127
transform 1 0 49518 0 1 130023
box -158 -213 158 213
use sky130_fd_pr__nfet_01v8_VT3ZQW  XM6_2
timestamp 1695667127
transform 1 0 49518 0 1 130493
box -158 -213 158 213
use sky130_fd_pr__nfet_01v8_VT3ZQW  XM6
timestamp 1695667127
transform 1 0 49518 0 1 129553
box -158 -213 158 213
use sky130_fd_pr__nfet_01v8_VT3ZQW  XM6_3
timestamp 1695667127
transform 1 0 49518 0 1 129083
box -158 -213 158 213
use sky130_fd_pr__pfet_01v8_7DHACV  XM7
timestamp 1695664993
transform 1 0 51712 0 1 26292
box -112 -9252 112 9252
use sky130_fd_pr__nfet_01v8_VT3ZQW  XM8_1
timestamp 1695667127
transform 1 0 49898 0 1 130023
box -158 -213 158 213
use sky130_fd_pr__nfet_01v8_VT3ZQW  XM8
timestamp 1695667127
transform 1 0 49898 0 1 130493
box -158 -213 158 213
use sky130_fd_pr__nfet_01v8_VT3ZQW  XM8_3
timestamp 1695667127
transform 1 0 49898 0 1 129083
box -158 -213 158 213
use sky130_fd_pr__pfet_01v8_F76D73  XM9_1
timestamp 1695663670
transform 1 0 99594 0 1 78822
box -1594 -61782 1594 61782
use sky130_fd_pr__pfet_01v8_F76D73  XM9_2
timestamp 1695663670
transform 1 0 85194 0 1 78822
box -1594 -61782 1594 61782
use sky130_fd_pr__pfet_01v8_F76D73  XM9_3
timestamp 1695663670
transform 1 0 77994 0 1 78822
box -1594 -61782 1594 61782
use sky130_fd_pr__pfet_01v8_F76D73  XM9_4
timestamp 1695663670
transform 1 0 92394 0 1 78822
box -1594 -61782 1594 61782
use sky130_fd_pr__pfet_01v8_E769TZ  XM9_dummy_1
timestamp 1695663670
transform 1 0 63594 0 1 78818
box -1594 -63018 1594 63018
use sky130_fd_pr__pfet_01v8_SLZ774  XM9_dummy_3
timestamp 1695663670
transform 1 0 67194 0 1 16400
box -1594 -600 1594 600
use sky130_fd_pr__pfet_01v8_ZLZ7XS  XM9_dummy_4
timestamp 1695663670
transform 1 0 70794 0 1 16400
box -1594 -600 1594 600
use sky130_fd_pr__pfet_01v8_ZLZ7XS  XM9_dummy_5
timestamp 1695663670
transform 1 0 74394 0 1 16400
box -1594 -600 1594 600
use sky130_fd_pr__pfet_01v8_ZLZ7XS  XM9_dummy_6
timestamp 1695663670
transform 1 0 77994 0 1 16400
box -1594 -600 1594 600
use sky130_fd_pr__pfet_01v8_ZLZ7XS  XM9_dummy_7
timestamp 1695663670
transform 1 0 81594 0 1 16400
box -1594 -600 1594 600
use sky130_fd_pr__pfet_01v8_ZLZ7XS  XM9_dummy_8
timestamp 1695663670
transform 1 0 85194 0 1 16400
box -1594 -600 1594 600
use sky130_fd_pr__pfet_01v8_ZLZ7XS  XM9_dummy_9
timestamp 1695663670
transform 1 0 88794 0 1 16400
box -1594 -600 1594 600
use sky130_fd_pr__pfet_01v8_ZLZ7XS  XM9_dummy_10
timestamp 1695663670
transform 1 0 92394 0 1 16400
box -1594 -600 1594 600
use sky130_fd_pr__pfet_01v8_ZLZ7XS  XM9_dummy_11
timestamp 1695663670
transform 1 0 95994 0 1 16400
box -1594 -600 1594 600
use sky130_fd_pr__pfet_01v8_ZLZ7XS  XM9_dummy_12
timestamp 1695663670
transform 1 0 99594 0 1 16400
box -1594 -600 1594 600
use sky130_fd_pr__pfet_01v8_ZLZ7XS  XM9_dummy_13
timestamp 1695663670
transform 1 0 74394 0 1 141240
box -1594 -600 1594 600
use sky130_fd_pr__pfet_01v8_ZLZ7XS  XM9_dummy_14
timestamp 1695663670
transform 1 0 85194 0 1 141240
box -1594 -600 1594 600
use sky130_fd_pr__pfet_01v8_ZLZ7XS  XM9_dummy_16
timestamp 1695663670
transform 1 0 77994 0 1 141240
box -1594 -600 1594 600
use sky130_fd_pr__pfet_01v8_ZLZ7XS  XM9_dummy_17
timestamp 1695663670
transform 1 0 67194 0 1 141240
box -1594 -600 1594 600
use sky130_fd_pr__pfet_01v8_ZLZ7XS  XM9_dummy_18
timestamp 1695663670
transform 1 0 88794 0 1 141240
box -1594 -600 1594 600
use sky130_fd_pr__pfet_01v8_ZLZ7XS  XM9_dummy_19
timestamp 1695663670
transform 1 0 81594 0 1 141240
box -1594 -600 1594 600
use sky130_fd_pr__pfet_01v8_ZLZ7XS  XM9_dummy_20
timestamp 1695663670
transform 1 0 92394 0 1 141240
box -1594 -600 1594 600
use sky130_fd_pr__pfet_01v8_ZLZ7XS  XM9_dummy_22
timestamp 1695663670
transform 1 0 95994 0 1 141240
box -1594 -600 1594 600
use sky130_fd_pr__pfet_01v8_F76D73  XM9
timestamp 1695663670
transform 1 0 70794 0 1 78822
box -1594 -61782 1594 61782
use sky130_fd_pr__pfet_01v8_ZLZ7XS  XM9_dummy_15
timestamp 1695663670
transform 1 0 70794 0 1 141240
box -1594 -600 1594 600
use sky130_fd_pr__pfet_01v8_UDM5A5  XM10
timestamp 1695665689
transform 1 0 45594 0 1 76892
box -594 -9252 594 9252
use sky130_fd_pr__nfet_01v8_QP5WRD  XM11
timestamp 1695666081
transform 1 0 49758 0 1 102334
box -558 -9114 558 9114
use sky130_fd_pr__nfet_01v8_QP5WRD  XM11_1
timestamp 1695666081
transform 1 0 45558 0 1 102334
box -558 -9114 558 9114
use sky130_fd_pr__pfet_01v8_RRU5GE  XM100_1
timestamp 1695665377
transform 1 0 49594 0 1 51076
box -394 -1836 394 1836
use sky130_fd_pr__pfet_01v8_P2UXFR  XM100_4
timestamp 1695665377
transform 1 0 48794 0 1 50458
box -394 -1218 394 1218
use sky130_fd_pr__pfet_01v8_RRUZAE  XM100_dummy_1
timestamp 1695665377
transform 1 0 46394 0 1 51072
box -394 -3072 394 3072
use sky130_fd_pr__pfet_01v8_P2UXFR  XM100_dummy_3
timestamp 1695665377
transform 1 0 47994 0 1 52938
box -394 -1218 394 1218
use sky130_fd_pr__pfet_01v8_P2UXFR  XM100_dummy_4
timestamp 1695665377
transform 1 0 48794 0 1 52938
box -394 -1218 394 1218
use sky130_fd_pr__pfet_01v8_C2U9V5  XM100_dummy_5
timestamp 1695665377
transform 1 0 47194 0 1 53550
box -394 -600 394 600
use sky130_fd_pr__pfet_01v8_C2U9V5  XM100_dummy_6
timestamp 1695665377
transform 1 0 49594 0 1 53560
box -394 -600 394 600
use sky130_fd_pr__pfet_01v8_C2U9V5  XM100_dummy_7
timestamp 1695665377
transform 1 0 48794 0 1 48600
box -394 -600 394 600
use sky130_fd_pr__pfet_01v8_C2U9V5  XM100_dummy_8
timestamp 1695665377
transform 1 0 47194 0 1 48600
box -394 -600 394 600
use sky130_fd_pr__pfet_01v8_C2U9V5  XM100_dummy_9
timestamp 1695665377
transform 1 0 47994 0 1 48600
box -394 -600 394 600
<< labels >>
flabel metal2 50928 130008 51126 130070 0 FreeSans 1600 0 0 0 bias21
flabel metal2 47172 129858 47470 130044 0 FreeSans 1600 0 0 0 bias3
flabel metal2 59050 142302 59318 142626 0 FreeSans 1600 0 0 0 bias1
flabel metal1 56686 65906 57592 66152 0 FreeSans 8000 0 0 0 m1m2
flabel metal1 48258 117074 48380 117368 0 FreeSans 8000 0 0 0 m3m4
flabel metal2 51774 65034 52322 65266 0 FreeSans 8000 0 0 0 m9m10
flabel metal1 51824 118482 51912 118858 0 FreeSans 8000 0 0 0 m11m12
flabel metal1 52140 35720 52180 35780 0 FreeSans 1600 0 0 0 dummy_5
flabel metal1 50720 47780 50760 47840 0 FreeSans 1600 0 0 0 dummy_100
flabel metal1 51740 67560 51780 67640 0 FreeSans 1600 0 0 0 dummy_2
flabel metal1 51720 93180 51780 93240 0 FreeSans 1600 0 0 0 dummy_3
flabel metal1 50800 130740 50820 130760 0 FreeSans 1600 0 0 0 dummy_4
flabel metal1 104760 16940 104820 17040 0 FreeSans 1600 0 0 0 dummy_9
flabel metal3 32800 112000 34800 114000 0 FreeSans 3200 0 0 0 VB_B
port 6 nsew signal bidirectional
flabel metal3 32800 90000 34800 92000 0 FreeSans 3200 0 0 0 OUT
port 4 nsew signal bidirectional
flabel metal3 32800 86000 34800 88000 0 FreeSans 3200 0 0 0 VB_A
port 5 nsew signal bidirectional
flabel metal3 32800 54000 34800 56000 0 FreeSans 3200 0 0 0 IB
port 7 nsew signal bidirectional
flabel metal3 32800 18000 34800 20000 0 FreeSans 3200 0 0 0 IN_M
port 1 nsew signal bidirectional
flabel metal3 32800 14000 34800 16000 0 FreeSans 3200 0 0 0 IN_P
port 0 nsew signal bidirectional
flabel metal3 32800 143000 34800 145000 0 FreeSans 3200 0 0 0 VSS
port 3 nsew ground bidirectional
flabel metal3 32800 139000 34800 141000 0 FreeSans 3200 0 0 0 VCC
port 2 nsew power bidirectional
<< end >>
